magic
tech scmos
timestamp 1638840038
<< nwell >>
rect 18 1377 74 1397
rect 117 1377 141 1397
rect 147 1377 203 1397
rect 238 1377 294 1397
rect 337 1377 361 1397
rect 367 1377 423 1397
rect 458 1377 514 1397
rect 557 1377 581 1397
rect 587 1377 643 1397
rect 678 1377 734 1397
rect 777 1377 801 1397
rect 807 1377 863 1397
rect 117 1327 141 1347
rect 337 1327 361 1347
rect 557 1327 581 1347
rect 777 1327 801 1347
rect 221 1115 277 1135
rect 331 1115 387 1135
rect 480 1115 536 1135
rect 670 1115 726 1135
rect 331 1052 399 1072
rect 480 1052 548 1072
rect 670 1052 738 1072
rect 480 982 560 1002
rect 670 982 750 1002
rect 670 905 762 925
rect 218 821 274 841
rect 328 821 396 841
rect 477 821 557 841
rect 667 821 759 841
rect 109 701 133 721
rect 139 701 195 721
rect 249 701 273 721
rect 279 701 335 721
rect 389 701 413 721
rect 419 701 475 721
rect 529 701 553 721
rect 559 701 615 721
rect 109 651 133 671
rect 249 651 273 671
rect 389 651 413 671
rect 529 651 553 671
<< ntransistor >>
rect 128 1365 130 1369
rect 31 1351 33 1355
rect 43 1351 45 1355
rect 61 1351 63 1355
rect 348 1365 350 1369
rect 251 1351 253 1355
rect 263 1351 265 1355
rect 281 1351 283 1355
rect 568 1365 570 1369
rect 471 1351 473 1355
rect 483 1351 485 1355
rect 501 1351 503 1355
rect 788 1365 790 1369
rect 691 1351 693 1355
rect 703 1351 705 1355
rect 721 1351 723 1355
rect 128 1315 130 1319
rect 159 1315 161 1319
rect 169 1315 171 1319
rect 179 1315 181 1319
rect 189 1315 191 1319
rect 348 1315 350 1319
rect 379 1315 381 1319
rect 389 1315 391 1319
rect 399 1315 401 1319
rect 409 1315 411 1319
rect 568 1315 570 1319
rect 599 1315 601 1319
rect 609 1315 611 1319
rect 619 1315 621 1319
rect 629 1315 631 1319
rect 788 1315 790 1319
rect 819 1315 821 1319
rect 829 1315 831 1319
rect 839 1315 841 1319
rect 849 1315 851 1319
rect 234 1089 236 1093
rect 246 1089 248 1093
rect 264 1089 266 1093
rect 344 1089 346 1093
rect 356 1089 358 1093
rect 374 1089 376 1093
rect 493 1089 495 1093
rect 505 1089 507 1093
rect 523 1089 525 1093
rect 683 1089 685 1093
rect 695 1089 697 1093
rect 713 1089 715 1093
rect 344 1019 346 1023
rect 356 1019 358 1023
rect 368 1019 370 1023
rect 386 1019 388 1023
rect 493 1019 495 1023
rect 505 1019 507 1023
rect 517 1019 519 1023
rect 535 1019 537 1023
rect 683 1019 685 1023
rect 695 1019 697 1023
rect 707 1019 709 1023
rect 725 1019 727 1023
rect 493 942 495 946
rect 505 942 507 946
rect 517 942 519 946
rect 529 942 531 946
rect 547 942 549 946
rect 683 942 685 946
rect 695 942 697 946
rect 707 942 709 946
rect 719 942 721 946
rect 737 942 739 946
rect 683 858 685 862
rect 695 858 697 862
rect 707 858 709 862
rect 719 858 721 862
rect 731 858 733 862
rect 749 858 751 862
rect 229 795 231 799
rect 247 795 249 799
rect 259 795 261 799
rect 339 788 341 792
rect 357 788 359 792
rect 369 788 371 792
rect 381 788 383 792
rect 488 781 490 785
rect 506 781 508 785
rect 518 781 520 785
rect 530 781 532 785
rect 542 781 544 785
rect 678 774 680 778
rect 696 774 698 778
rect 708 774 710 778
rect 720 774 722 778
rect 732 774 734 778
rect 744 774 746 778
rect 120 689 122 693
rect 260 689 262 693
rect 400 689 402 693
rect 540 689 542 693
rect 120 639 122 643
rect 151 639 153 643
rect 161 639 163 643
rect 171 639 173 643
rect 181 639 183 643
rect 260 639 262 643
rect 291 639 293 643
rect 301 639 303 643
rect 311 639 313 643
rect 321 639 323 643
rect 400 639 402 643
rect 431 639 433 643
rect 441 639 443 643
rect 451 639 453 643
rect 461 639 463 643
rect 540 639 542 643
rect 571 639 573 643
rect 581 639 583 643
rect 591 639 593 643
rect 601 639 603 643
<< ptransistor >>
rect 31 1383 33 1391
rect 43 1383 45 1391
rect 61 1383 63 1391
rect 128 1383 130 1391
rect 159 1383 161 1391
rect 169 1383 171 1391
rect 179 1383 181 1391
rect 189 1383 191 1391
rect 128 1333 130 1341
rect 251 1383 253 1391
rect 263 1383 265 1391
rect 281 1383 283 1391
rect 348 1383 350 1391
rect 379 1383 381 1391
rect 389 1383 391 1391
rect 399 1383 401 1391
rect 409 1383 411 1391
rect 348 1333 350 1341
rect 471 1383 473 1391
rect 483 1383 485 1391
rect 501 1383 503 1391
rect 568 1383 570 1391
rect 599 1383 601 1391
rect 609 1383 611 1391
rect 619 1383 621 1391
rect 629 1383 631 1391
rect 568 1333 570 1341
rect 691 1383 693 1391
rect 703 1383 705 1391
rect 721 1383 723 1391
rect 788 1383 790 1391
rect 819 1383 821 1391
rect 829 1383 831 1391
rect 839 1383 841 1391
rect 849 1383 851 1391
rect 788 1333 790 1341
rect 234 1121 236 1129
rect 246 1121 248 1129
rect 264 1121 266 1129
rect 344 1121 346 1129
rect 356 1121 358 1129
rect 374 1121 376 1129
rect 493 1121 495 1129
rect 505 1121 507 1129
rect 523 1121 525 1129
rect 683 1121 685 1129
rect 695 1121 697 1129
rect 713 1121 715 1129
rect 344 1058 346 1066
rect 356 1058 358 1066
rect 368 1058 370 1066
rect 386 1058 388 1066
rect 493 1058 495 1066
rect 505 1058 507 1066
rect 517 1058 519 1066
rect 535 1058 537 1066
rect 683 1058 685 1066
rect 695 1058 697 1066
rect 707 1058 709 1066
rect 725 1058 727 1066
rect 493 988 495 996
rect 505 988 507 996
rect 517 988 519 996
rect 529 988 531 996
rect 547 988 549 996
rect 683 988 685 996
rect 695 988 697 996
rect 707 988 709 996
rect 719 988 721 996
rect 737 988 739 996
rect 683 911 685 919
rect 695 911 697 919
rect 707 911 709 919
rect 719 911 721 919
rect 731 911 733 919
rect 749 911 751 919
rect 229 827 231 835
rect 247 827 249 835
rect 259 827 261 835
rect 339 827 341 835
rect 357 827 359 835
rect 369 827 371 835
rect 381 827 383 835
rect 488 827 490 835
rect 506 827 508 835
rect 518 827 520 835
rect 530 827 532 835
rect 542 827 544 835
rect 678 827 680 835
rect 696 827 698 835
rect 708 827 710 835
rect 720 827 722 835
rect 732 827 734 835
rect 744 827 746 835
rect 120 707 122 715
rect 151 707 153 715
rect 161 707 163 715
rect 171 707 173 715
rect 181 707 183 715
rect 120 657 122 665
rect 260 707 262 715
rect 291 707 293 715
rect 301 707 303 715
rect 311 707 313 715
rect 321 707 323 715
rect 260 657 262 665
rect 400 707 402 715
rect 431 707 433 715
rect 441 707 443 715
rect 451 707 453 715
rect 461 707 463 715
rect 400 657 402 665
rect 540 707 542 715
rect 571 707 573 715
rect 581 707 583 715
rect 591 707 593 715
rect 601 707 603 715
rect 540 657 542 665
<< ndiffusion >>
rect 127 1365 128 1369
rect 130 1365 131 1369
rect 28 1351 31 1355
rect 33 1351 43 1355
rect 45 1351 48 1355
rect 60 1351 61 1355
rect 63 1351 64 1355
rect 347 1365 348 1369
rect 350 1365 351 1369
rect 248 1351 251 1355
rect 253 1351 263 1355
rect 265 1351 268 1355
rect 280 1351 281 1355
rect 283 1351 284 1355
rect 567 1365 568 1369
rect 570 1365 571 1369
rect 468 1351 471 1355
rect 473 1351 483 1355
rect 485 1351 488 1355
rect 500 1351 501 1355
rect 503 1351 504 1355
rect 787 1365 788 1369
rect 790 1365 791 1369
rect 688 1351 691 1355
rect 693 1351 703 1355
rect 705 1351 708 1355
rect 720 1351 721 1355
rect 723 1351 724 1355
rect 127 1315 128 1319
rect 130 1315 131 1319
rect 157 1315 159 1319
rect 161 1315 169 1319
rect 171 1315 173 1319
rect 177 1315 179 1319
rect 181 1315 189 1319
rect 191 1315 193 1319
rect 347 1315 348 1319
rect 350 1315 351 1319
rect 377 1315 379 1319
rect 381 1315 389 1319
rect 391 1315 393 1319
rect 397 1315 399 1319
rect 401 1315 409 1319
rect 411 1315 413 1319
rect 567 1315 568 1319
rect 570 1315 571 1319
rect 597 1315 599 1319
rect 601 1315 609 1319
rect 611 1315 613 1319
rect 617 1315 619 1319
rect 621 1315 629 1319
rect 631 1315 633 1319
rect 787 1315 788 1319
rect 790 1315 791 1319
rect 817 1315 819 1319
rect 821 1315 829 1319
rect 831 1315 833 1319
rect 837 1315 839 1319
rect 841 1315 849 1319
rect 851 1315 853 1319
rect 231 1089 234 1093
rect 236 1089 246 1093
rect 248 1089 251 1093
rect 263 1089 264 1093
rect 266 1089 267 1093
rect 341 1089 344 1093
rect 346 1089 356 1093
rect 358 1089 361 1093
rect 373 1089 374 1093
rect 376 1089 377 1093
rect 490 1089 493 1093
rect 495 1089 505 1093
rect 507 1089 510 1093
rect 522 1089 523 1093
rect 525 1089 526 1093
rect 680 1089 683 1093
rect 685 1089 695 1093
rect 697 1089 700 1093
rect 712 1089 713 1093
rect 715 1089 716 1093
rect 341 1019 344 1023
rect 346 1019 356 1023
rect 358 1019 368 1023
rect 370 1019 373 1023
rect 385 1019 386 1023
rect 388 1019 389 1023
rect 490 1019 493 1023
rect 495 1019 505 1023
rect 507 1019 517 1023
rect 519 1019 522 1023
rect 534 1019 535 1023
rect 537 1019 538 1023
rect 680 1019 683 1023
rect 685 1019 695 1023
rect 697 1019 707 1023
rect 709 1019 712 1023
rect 724 1019 725 1023
rect 727 1019 728 1023
rect 490 942 493 946
rect 495 942 505 946
rect 507 942 517 946
rect 519 942 529 946
rect 531 942 534 946
rect 546 942 547 946
rect 549 942 550 946
rect 680 942 683 946
rect 685 942 695 946
rect 697 942 707 946
rect 709 942 719 946
rect 721 942 724 946
rect 736 942 737 946
rect 739 942 740 946
rect 680 858 683 862
rect 685 858 695 862
rect 697 858 707 862
rect 709 858 719 862
rect 721 858 731 862
rect 733 858 736 862
rect 748 858 749 862
rect 751 858 752 862
rect 228 795 229 799
rect 231 795 232 799
rect 244 795 247 799
rect 249 795 252 799
rect 256 795 259 799
rect 261 795 264 799
rect 338 788 339 792
rect 341 788 342 792
rect 354 788 357 792
rect 359 788 362 792
rect 366 788 369 792
rect 371 788 374 792
rect 378 788 381 792
rect 383 788 386 792
rect 487 781 488 785
rect 490 781 491 785
rect 503 781 506 785
rect 508 781 511 785
rect 515 781 518 785
rect 520 781 523 785
rect 527 781 530 785
rect 532 781 535 785
rect 539 781 542 785
rect 544 781 547 785
rect 677 774 678 778
rect 680 774 681 778
rect 693 774 696 778
rect 698 774 701 778
rect 705 774 708 778
rect 710 774 713 778
rect 717 774 720 778
rect 722 774 725 778
rect 729 774 732 778
rect 734 774 737 778
rect 741 774 744 778
rect 746 774 749 778
rect 119 689 120 693
rect 122 689 123 693
rect 259 689 260 693
rect 262 689 263 693
rect 399 689 400 693
rect 402 689 403 693
rect 539 689 540 693
rect 542 689 543 693
rect 119 639 120 643
rect 122 639 123 643
rect 149 639 151 643
rect 153 639 161 643
rect 163 639 165 643
rect 169 639 171 643
rect 173 639 181 643
rect 183 639 185 643
rect 259 639 260 643
rect 262 639 263 643
rect 289 639 291 643
rect 293 639 301 643
rect 303 639 305 643
rect 309 639 311 643
rect 313 639 321 643
rect 323 639 325 643
rect 399 639 400 643
rect 402 639 403 643
rect 429 639 431 643
rect 433 639 441 643
rect 443 639 445 643
rect 449 639 451 643
rect 453 639 461 643
rect 463 639 465 643
rect 539 639 540 643
rect 542 639 543 643
rect 569 639 571 643
rect 573 639 581 643
rect 583 639 585 643
rect 589 639 591 643
rect 593 639 601 643
rect 603 639 605 643
<< pdiffusion >>
rect 28 1383 31 1391
rect 33 1383 36 1391
rect 40 1383 43 1391
rect 45 1383 48 1391
rect 60 1383 61 1391
rect 63 1383 64 1391
rect 127 1383 128 1391
rect 130 1383 131 1391
rect 157 1383 159 1391
rect 161 1383 169 1391
rect 171 1383 173 1391
rect 177 1383 179 1391
rect 181 1383 189 1391
rect 191 1383 193 1391
rect 127 1333 128 1341
rect 130 1333 131 1341
rect 248 1383 251 1391
rect 253 1383 256 1391
rect 260 1383 263 1391
rect 265 1383 268 1391
rect 280 1383 281 1391
rect 283 1383 284 1391
rect 347 1383 348 1391
rect 350 1383 351 1391
rect 377 1383 379 1391
rect 381 1383 389 1391
rect 391 1383 393 1391
rect 397 1383 399 1391
rect 401 1383 409 1391
rect 411 1383 413 1391
rect 347 1333 348 1341
rect 350 1333 351 1341
rect 468 1383 471 1391
rect 473 1383 476 1391
rect 480 1383 483 1391
rect 485 1383 488 1391
rect 500 1383 501 1391
rect 503 1383 504 1391
rect 567 1383 568 1391
rect 570 1383 571 1391
rect 597 1383 599 1391
rect 601 1383 609 1391
rect 611 1383 613 1391
rect 617 1383 619 1391
rect 621 1383 629 1391
rect 631 1383 633 1391
rect 567 1333 568 1341
rect 570 1333 571 1341
rect 688 1383 691 1391
rect 693 1383 696 1391
rect 700 1383 703 1391
rect 705 1383 708 1391
rect 720 1383 721 1391
rect 723 1383 724 1391
rect 787 1383 788 1391
rect 790 1383 791 1391
rect 817 1383 819 1391
rect 821 1383 829 1391
rect 831 1383 833 1391
rect 837 1383 839 1391
rect 841 1383 849 1391
rect 851 1383 853 1391
rect 787 1333 788 1341
rect 790 1333 791 1341
rect 231 1121 234 1129
rect 236 1121 239 1129
rect 243 1121 246 1129
rect 248 1121 251 1129
rect 263 1121 264 1129
rect 266 1121 267 1129
rect 341 1121 344 1129
rect 346 1121 349 1129
rect 353 1121 356 1129
rect 358 1121 361 1129
rect 373 1121 374 1129
rect 376 1121 377 1129
rect 490 1121 493 1129
rect 495 1121 498 1129
rect 502 1121 505 1129
rect 507 1121 510 1129
rect 522 1121 523 1129
rect 525 1121 526 1129
rect 680 1121 683 1129
rect 685 1121 688 1129
rect 692 1121 695 1129
rect 697 1121 700 1129
rect 712 1121 713 1129
rect 715 1121 716 1129
rect 341 1058 344 1066
rect 346 1058 349 1066
rect 353 1058 356 1066
rect 358 1058 361 1066
rect 365 1058 368 1066
rect 370 1058 373 1066
rect 385 1058 386 1066
rect 388 1058 389 1066
rect 490 1058 493 1066
rect 495 1058 498 1066
rect 502 1058 505 1066
rect 507 1058 510 1066
rect 514 1058 517 1066
rect 519 1058 522 1066
rect 534 1058 535 1066
rect 537 1058 538 1066
rect 680 1058 683 1066
rect 685 1058 688 1066
rect 692 1058 695 1066
rect 697 1058 700 1066
rect 704 1058 707 1066
rect 709 1058 712 1066
rect 724 1058 725 1066
rect 727 1058 728 1066
rect 490 988 493 996
rect 495 988 498 996
rect 502 988 505 996
rect 507 988 510 996
rect 514 988 517 996
rect 519 988 522 996
rect 526 988 529 996
rect 531 988 534 996
rect 546 988 547 996
rect 549 988 550 996
rect 680 988 683 996
rect 685 988 688 996
rect 692 988 695 996
rect 697 988 700 996
rect 704 988 707 996
rect 709 988 712 996
rect 716 988 719 996
rect 721 988 724 996
rect 736 988 737 996
rect 739 988 740 996
rect 680 911 683 919
rect 685 911 688 919
rect 692 911 695 919
rect 697 911 700 919
rect 704 911 707 919
rect 709 911 712 919
rect 716 911 719 919
rect 721 911 724 919
rect 728 911 731 919
rect 733 911 736 919
rect 748 911 749 919
rect 751 911 752 919
rect 228 827 229 835
rect 231 827 232 835
rect 244 827 247 835
rect 249 827 259 835
rect 261 827 264 835
rect 338 827 339 835
rect 341 827 342 835
rect 354 827 357 835
rect 359 827 369 835
rect 371 827 381 835
rect 383 827 386 835
rect 487 827 488 835
rect 490 827 491 835
rect 503 827 506 835
rect 508 827 518 835
rect 520 827 530 835
rect 532 827 542 835
rect 544 827 547 835
rect 677 827 678 835
rect 680 827 681 835
rect 693 827 696 835
rect 698 827 708 835
rect 710 827 720 835
rect 722 827 732 835
rect 734 827 744 835
rect 746 827 749 835
rect 119 707 120 715
rect 122 707 123 715
rect 149 707 151 715
rect 153 707 161 715
rect 163 707 165 715
rect 169 707 171 715
rect 173 707 181 715
rect 183 707 185 715
rect 119 657 120 665
rect 122 657 123 665
rect 259 707 260 715
rect 262 707 263 715
rect 289 707 291 715
rect 293 707 301 715
rect 303 707 305 715
rect 309 707 311 715
rect 313 707 321 715
rect 323 707 325 715
rect 259 657 260 665
rect 262 657 263 665
rect 399 707 400 715
rect 402 707 403 715
rect 429 707 431 715
rect 433 707 441 715
rect 443 707 445 715
rect 449 707 451 715
rect 453 707 461 715
rect 463 707 465 715
rect 399 657 400 665
rect 402 657 403 665
rect 539 707 540 715
rect 542 707 543 715
rect 569 707 571 715
rect 573 707 581 715
rect 583 707 585 715
rect 589 707 591 715
rect 593 707 601 715
rect 603 707 605 715
rect 539 657 540 665
rect 542 657 543 665
<< ndcontact >>
rect 123 1365 127 1369
rect 131 1365 135 1369
rect 24 1351 28 1355
rect 48 1351 52 1355
rect 56 1351 60 1355
rect 64 1351 68 1355
rect 343 1365 347 1369
rect 351 1365 355 1369
rect 244 1351 248 1355
rect 268 1351 272 1355
rect 276 1351 280 1355
rect 284 1351 288 1355
rect 563 1365 567 1369
rect 571 1365 575 1369
rect 464 1351 468 1355
rect 488 1351 492 1355
rect 496 1351 500 1355
rect 504 1351 508 1355
rect 783 1365 787 1369
rect 791 1365 795 1369
rect 684 1351 688 1355
rect 708 1351 712 1355
rect 716 1351 720 1355
rect 724 1351 728 1355
rect 123 1315 127 1319
rect 131 1315 135 1319
rect 153 1315 157 1319
rect 173 1315 177 1319
rect 193 1315 197 1319
rect 343 1315 347 1319
rect 351 1315 355 1319
rect 373 1315 377 1319
rect 393 1315 397 1319
rect 413 1315 417 1319
rect 563 1315 567 1319
rect 571 1315 575 1319
rect 593 1315 597 1319
rect 613 1315 617 1319
rect 633 1315 637 1319
rect 783 1315 787 1319
rect 791 1315 795 1319
rect 813 1315 817 1319
rect 833 1315 837 1319
rect 853 1315 857 1319
rect 227 1089 231 1093
rect 251 1089 255 1093
rect 259 1089 263 1093
rect 267 1089 271 1093
rect 337 1089 341 1093
rect 361 1089 365 1093
rect 369 1089 373 1093
rect 377 1089 381 1093
rect 486 1089 490 1093
rect 510 1089 514 1093
rect 518 1089 522 1093
rect 526 1089 530 1093
rect 676 1089 680 1093
rect 700 1089 704 1093
rect 708 1089 712 1093
rect 716 1089 720 1093
rect 337 1019 341 1023
rect 373 1019 377 1023
rect 381 1019 385 1023
rect 389 1019 393 1023
rect 486 1019 490 1023
rect 522 1019 526 1023
rect 530 1019 534 1023
rect 538 1019 542 1023
rect 676 1019 680 1023
rect 712 1019 716 1023
rect 720 1019 724 1023
rect 728 1019 732 1023
rect 486 942 490 946
rect 534 942 538 946
rect 542 942 546 946
rect 550 942 554 946
rect 676 942 680 946
rect 724 942 728 946
rect 732 942 736 946
rect 740 942 744 946
rect 676 858 680 862
rect 736 858 740 862
rect 744 858 748 862
rect 752 858 756 862
rect 224 795 228 799
rect 232 795 236 799
rect 240 795 244 799
rect 252 795 256 799
rect 264 795 268 799
rect 334 788 338 792
rect 342 788 346 792
rect 350 788 354 792
rect 362 788 366 792
rect 374 788 378 792
rect 386 788 390 792
rect 483 781 487 785
rect 491 781 495 785
rect 499 781 503 785
rect 511 781 515 785
rect 523 781 527 785
rect 535 781 539 785
rect 547 781 551 785
rect 673 774 677 778
rect 681 774 685 778
rect 689 774 693 778
rect 701 774 705 778
rect 713 774 717 778
rect 725 774 729 778
rect 737 774 741 778
rect 749 774 753 778
rect 115 689 119 693
rect 123 689 127 693
rect 255 689 259 693
rect 263 689 267 693
rect 395 689 399 693
rect 403 689 407 693
rect 535 689 539 693
rect 543 689 547 693
rect 115 639 119 643
rect 123 639 127 643
rect 145 639 149 643
rect 165 639 169 643
rect 185 639 189 643
rect 255 639 259 643
rect 263 639 267 643
rect 285 639 289 643
rect 305 639 309 643
rect 325 639 329 643
rect 395 639 399 643
rect 403 639 407 643
rect 425 639 429 643
rect 445 639 449 643
rect 465 639 469 643
rect 535 639 539 643
rect 543 639 547 643
rect 565 639 569 643
rect 585 639 589 643
rect 605 639 609 643
<< pdcontact >>
rect 24 1383 28 1391
rect 36 1383 40 1391
rect 48 1383 52 1391
rect 56 1383 60 1391
rect 64 1383 68 1391
rect 123 1383 127 1391
rect 131 1383 135 1391
rect 153 1383 157 1391
rect 173 1383 177 1391
rect 193 1383 197 1391
rect 123 1333 127 1341
rect 131 1333 135 1341
rect 244 1383 248 1391
rect 256 1383 260 1391
rect 268 1383 272 1391
rect 276 1383 280 1391
rect 284 1383 288 1391
rect 343 1383 347 1391
rect 351 1383 355 1391
rect 373 1383 377 1391
rect 393 1383 397 1391
rect 413 1383 417 1391
rect 343 1333 347 1341
rect 351 1333 355 1341
rect 464 1383 468 1391
rect 476 1383 480 1391
rect 488 1383 492 1391
rect 496 1383 500 1391
rect 504 1383 508 1391
rect 563 1383 567 1391
rect 571 1383 575 1391
rect 593 1383 597 1391
rect 613 1383 617 1391
rect 633 1383 637 1391
rect 563 1333 567 1341
rect 571 1333 575 1341
rect 684 1383 688 1391
rect 696 1383 700 1391
rect 708 1383 712 1391
rect 716 1383 720 1391
rect 724 1383 728 1391
rect 783 1383 787 1391
rect 791 1383 795 1391
rect 813 1383 817 1391
rect 833 1383 837 1391
rect 853 1383 857 1391
rect 783 1333 787 1341
rect 791 1333 795 1341
rect 227 1121 231 1129
rect 239 1121 243 1129
rect 251 1121 255 1129
rect 259 1121 263 1129
rect 267 1121 271 1129
rect 337 1121 341 1129
rect 349 1121 353 1129
rect 361 1121 365 1129
rect 369 1121 373 1129
rect 377 1121 381 1129
rect 486 1121 490 1129
rect 498 1121 502 1129
rect 510 1121 514 1129
rect 518 1121 522 1129
rect 526 1121 530 1129
rect 676 1121 680 1129
rect 688 1121 692 1129
rect 700 1121 704 1129
rect 708 1121 712 1129
rect 716 1121 720 1129
rect 337 1058 341 1066
rect 349 1058 353 1066
rect 361 1058 365 1066
rect 373 1058 377 1066
rect 381 1058 385 1066
rect 389 1058 393 1066
rect 486 1058 490 1066
rect 498 1058 502 1066
rect 510 1058 514 1066
rect 522 1058 526 1066
rect 530 1058 534 1066
rect 538 1058 542 1066
rect 676 1058 680 1066
rect 688 1058 692 1066
rect 700 1058 704 1066
rect 712 1058 716 1066
rect 720 1058 724 1066
rect 728 1058 732 1066
rect 486 988 490 996
rect 498 988 502 996
rect 510 988 514 996
rect 522 988 526 996
rect 534 988 538 996
rect 542 988 546 996
rect 550 988 554 996
rect 676 988 680 996
rect 688 988 692 996
rect 700 988 704 996
rect 712 988 716 996
rect 724 988 728 996
rect 732 988 736 996
rect 740 988 744 996
rect 676 911 680 919
rect 688 911 692 919
rect 700 911 704 919
rect 712 911 716 919
rect 724 911 728 919
rect 736 911 740 919
rect 744 911 748 919
rect 752 911 756 919
rect 224 827 228 835
rect 232 827 236 835
rect 240 827 244 835
rect 264 827 268 835
rect 334 827 338 835
rect 342 827 346 835
rect 350 827 354 835
rect 386 827 390 835
rect 483 827 487 835
rect 491 827 495 835
rect 499 827 503 835
rect 547 827 551 835
rect 673 827 677 835
rect 681 827 685 835
rect 689 827 693 835
rect 749 827 753 835
rect 115 707 119 715
rect 123 707 127 715
rect 145 707 149 715
rect 165 707 169 715
rect 185 707 189 715
rect 115 657 119 665
rect 123 657 127 665
rect 255 707 259 715
rect 263 707 267 715
rect 285 707 289 715
rect 305 707 309 715
rect 325 707 329 715
rect 255 657 259 665
rect 263 657 267 665
rect 395 707 399 715
rect 403 707 407 715
rect 425 707 429 715
rect 445 707 449 715
rect 465 707 469 715
rect 395 657 399 665
rect 403 657 407 665
rect 535 707 539 715
rect 543 707 547 715
rect 565 707 569 715
rect 585 707 589 715
rect 605 707 609 715
rect 535 657 539 665
rect 543 657 547 665
<< polysilicon >>
rect 159 1401 201 1403
rect 31 1391 33 1394
rect 43 1391 45 1394
rect 61 1391 63 1394
rect 128 1391 130 1394
rect 159 1391 161 1401
rect 169 1391 171 1394
rect 179 1391 181 1394
rect 189 1391 191 1394
rect 31 1355 33 1383
rect 43 1355 45 1383
rect 61 1355 63 1383
rect 128 1369 130 1383
rect 159 1372 161 1383
rect 169 1368 171 1383
rect 159 1366 171 1368
rect 128 1362 130 1365
rect 31 1348 33 1351
rect 43 1348 45 1351
rect 61 1348 63 1351
rect 128 1341 130 1344
rect 128 1319 130 1333
rect 159 1319 161 1366
rect 179 1363 181 1383
rect 169 1361 181 1363
rect 169 1319 171 1361
rect 189 1329 191 1383
rect 179 1327 191 1329
rect 179 1319 181 1327
rect 199 1324 201 1401
rect 379 1401 421 1403
rect 251 1391 253 1394
rect 263 1391 265 1394
rect 281 1391 283 1394
rect 348 1391 350 1394
rect 379 1391 381 1401
rect 389 1391 391 1394
rect 399 1391 401 1394
rect 409 1391 411 1394
rect 251 1355 253 1383
rect 263 1355 265 1383
rect 281 1355 283 1383
rect 348 1369 350 1383
rect 379 1372 381 1383
rect 389 1368 391 1383
rect 379 1366 391 1368
rect 348 1362 350 1365
rect 251 1348 253 1351
rect 263 1348 265 1351
rect 281 1348 283 1351
rect 348 1341 350 1344
rect 189 1322 201 1324
rect 189 1319 191 1322
rect 348 1319 350 1333
rect 379 1319 381 1366
rect 399 1363 401 1383
rect 389 1361 401 1363
rect 389 1319 391 1361
rect 409 1329 411 1383
rect 399 1327 411 1329
rect 399 1319 401 1327
rect 419 1324 421 1401
rect 599 1401 641 1403
rect 471 1391 473 1394
rect 483 1391 485 1394
rect 501 1391 503 1394
rect 568 1391 570 1394
rect 599 1391 601 1401
rect 609 1391 611 1394
rect 619 1391 621 1394
rect 629 1391 631 1394
rect 471 1355 473 1383
rect 483 1355 485 1383
rect 501 1355 503 1383
rect 568 1369 570 1383
rect 599 1372 601 1383
rect 609 1368 611 1383
rect 599 1366 611 1368
rect 568 1362 570 1365
rect 471 1348 473 1351
rect 483 1348 485 1351
rect 501 1348 503 1351
rect 568 1341 570 1344
rect 409 1322 421 1324
rect 409 1319 411 1322
rect 568 1319 570 1333
rect 599 1319 601 1366
rect 619 1363 621 1383
rect 609 1361 621 1363
rect 609 1319 611 1361
rect 629 1329 631 1383
rect 619 1327 631 1329
rect 619 1319 621 1327
rect 639 1324 641 1401
rect 819 1401 861 1403
rect 691 1391 693 1394
rect 703 1391 705 1394
rect 721 1391 723 1394
rect 788 1391 790 1394
rect 819 1391 821 1401
rect 829 1391 831 1394
rect 839 1391 841 1394
rect 849 1391 851 1394
rect 691 1355 693 1383
rect 703 1355 705 1383
rect 721 1355 723 1383
rect 788 1369 790 1383
rect 819 1372 821 1383
rect 829 1368 831 1383
rect 819 1366 831 1368
rect 788 1362 790 1365
rect 691 1348 693 1351
rect 703 1348 705 1351
rect 721 1348 723 1351
rect 788 1341 790 1344
rect 629 1322 641 1324
rect 629 1319 631 1322
rect 788 1319 790 1333
rect 819 1319 821 1366
rect 839 1363 841 1383
rect 829 1361 841 1363
rect 829 1319 831 1361
rect 849 1329 851 1383
rect 839 1327 851 1329
rect 839 1319 841 1327
rect 859 1324 861 1401
rect 849 1322 861 1324
rect 849 1319 851 1322
rect 128 1312 130 1315
rect 159 1299 161 1315
rect 169 1312 171 1315
rect 179 1291 181 1315
rect 189 1312 191 1315
rect 348 1312 350 1315
rect 379 1299 381 1315
rect 389 1312 391 1315
rect 399 1291 401 1315
rect 409 1312 411 1315
rect 568 1312 570 1315
rect 599 1299 601 1315
rect 609 1312 611 1315
rect 619 1291 621 1315
rect 629 1312 631 1315
rect 788 1312 790 1315
rect 819 1299 821 1315
rect 829 1312 831 1315
rect 839 1291 841 1315
rect 849 1312 851 1315
rect 234 1129 236 1132
rect 246 1129 248 1132
rect 264 1129 266 1132
rect 344 1129 346 1132
rect 356 1129 358 1132
rect 374 1129 376 1132
rect 493 1129 495 1132
rect 505 1129 507 1132
rect 523 1129 525 1132
rect 683 1129 685 1132
rect 695 1129 697 1132
rect 713 1129 715 1132
rect 234 1093 236 1121
rect 246 1093 248 1121
rect 264 1093 266 1121
rect 344 1093 346 1121
rect 356 1093 358 1121
rect 374 1093 376 1121
rect 493 1093 495 1121
rect 505 1093 507 1121
rect 523 1093 525 1121
rect 683 1093 685 1121
rect 695 1093 697 1121
rect 713 1093 715 1121
rect 234 1086 236 1089
rect 246 1086 248 1089
rect 264 1086 266 1089
rect 344 1086 346 1089
rect 356 1086 358 1089
rect 374 1086 376 1089
rect 493 1086 495 1089
rect 505 1086 507 1089
rect 523 1086 525 1089
rect 683 1086 685 1089
rect 695 1086 697 1089
rect 713 1086 715 1089
rect 344 1066 346 1069
rect 356 1066 358 1069
rect 368 1066 370 1069
rect 386 1066 388 1069
rect 493 1066 495 1069
rect 505 1066 507 1069
rect 517 1066 519 1069
rect 535 1066 537 1069
rect 683 1066 685 1069
rect 695 1066 697 1069
rect 707 1066 709 1069
rect 725 1066 727 1069
rect 344 1023 346 1058
rect 356 1023 358 1058
rect 368 1023 370 1058
rect 386 1023 388 1058
rect 493 1023 495 1058
rect 505 1023 507 1058
rect 517 1023 519 1058
rect 535 1023 537 1058
rect 683 1023 685 1058
rect 695 1023 697 1058
rect 707 1023 709 1058
rect 725 1023 727 1058
rect 344 1016 346 1019
rect 356 1016 358 1019
rect 368 1016 370 1019
rect 386 1016 388 1019
rect 493 1016 495 1019
rect 505 1016 507 1019
rect 517 1016 519 1019
rect 535 1016 537 1019
rect 683 1016 685 1019
rect 695 1016 697 1019
rect 707 1016 709 1019
rect 725 1016 727 1019
rect 493 996 495 999
rect 505 996 507 999
rect 517 996 519 999
rect 529 996 531 999
rect 547 996 549 999
rect 683 996 685 999
rect 695 996 697 999
rect 707 996 709 999
rect 719 996 721 999
rect 737 996 739 999
rect 493 946 495 988
rect 505 946 507 988
rect 517 946 519 988
rect 529 946 531 988
rect 547 946 549 988
rect 683 946 685 988
rect 695 946 697 988
rect 707 946 709 988
rect 719 946 721 988
rect 737 946 739 988
rect 493 939 495 942
rect 505 939 507 942
rect 517 939 519 942
rect 529 939 531 942
rect 547 939 549 942
rect 683 939 685 942
rect 695 939 697 942
rect 707 939 709 942
rect 719 939 721 942
rect 737 939 739 942
rect 683 919 685 922
rect 695 919 697 922
rect 707 919 709 922
rect 719 919 721 922
rect 731 919 733 922
rect 749 919 751 922
rect 683 862 685 911
rect 695 862 697 911
rect 707 862 709 911
rect 719 862 721 911
rect 731 862 733 911
rect 749 862 751 911
rect 683 855 685 858
rect 695 855 697 858
rect 707 855 709 858
rect 719 855 721 858
rect 731 855 733 858
rect 749 855 751 858
rect 229 835 231 838
rect 247 835 249 838
rect 259 835 261 838
rect 339 835 341 838
rect 357 835 359 838
rect 369 835 371 838
rect 381 835 383 838
rect 488 835 490 838
rect 506 835 508 838
rect 518 835 520 838
rect 530 835 532 838
rect 542 835 544 838
rect 678 835 680 838
rect 696 835 698 838
rect 708 835 710 838
rect 720 835 722 838
rect 732 835 734 838
rect 744 835 746 838
rect 229 799 231 827
rect 247 799 249 827
rect 259 799 261 827
rect 229 792 231 795
rect 247 792 249 795
rect 259 792 261 795
rect 339 792 341 827
rect 357 792 359 827
rect 369 792 371 827
rect 381 792 383 827
rect 339 785 341 788
rect 357 785 359 788
rect 369 785 371 788
rect 381 785 383 788
rect 488 785 490 827
rect 506 785 508 827
rect 518 785 520 827
rect 530 785 532 827
rect 542 785 544 827
rect 488 778 490 781
rect 506 778 508 781
rect 518 778 520 781
rect 530 778 532 781
rect 542 778 544 781
rect 678 778 680 827
rect 696 778 698 827
rect 708 778 710 827
rect 720 778 722 827
rect 732 778 734 827
rect 744 778 746 827
rect 678 771 680 774
rect 696 771 698 774
rect 708 771 710 774
rect 720 771 722 774
rect 732 771 734 774
rect 744 771 746 774
rect 151 725 193 727
rect 120 715 122 718
rect 151 715 153 725
rect 161 715 163 718
rect 171 715 173 718
rect 181 715 183 718
rect 120 693 122 707
rect 151 696 153 707
rect 161 692 163 707
rect 151 690 163 692
rect 120 686 122 689
rect 120 665 122 668
rect 120 643 122 657
rect 151 643 153 690
rect 171 687 173 707
rect 161 685 173 687
rect 161 643 163 685
rect 181 653 183 707
rect 171 651 183 653
rect 171 643 173 651
rect 191 648 193 725
rect 291 725 333 727
rect 260 715 262 718
rect 291 715 293 725
rect 301 715 303 718
rect 311 715 313 718
rect 321 715 323 718
rect 260 693 262 707
rect 291 696 293 707
rect 301 692 303 707
rect 291 690 303 692
rect 260 686 262 689
rect 260 665 262 668
rect 181 646 193 648
rect 181 643 183 646
rect 260 643 262 657
rect 291 643 293 690
rect 311 687 313 707
rect 301 685 313 687
rect 301 643 303 685
rect 321 653 323 707
rect 311 651 323 653
rect 311 643 313 651
rect 331 648 333 725
rect 431 725 473 727
rect 400 715 402 718
rect 431 715 433 725
rect 441 715 443 718
rect 451 715 453 718
rect 461 715 463 718
rect 400 693 402 707
rect 431 696 433 707
rect 441 692 443 707
rect 431 690 443 692
rect 400 686 402 689
rect 400 665 402 668
rect 321 646 333 648
rect 321 643 323 646
rect 400 643 402 657
rect 431 643 433 690
rect 451 687 453 707
rect 441 685 453 687
rect 441 643 443 685
rect 461 653 463 707
rect 451 651 463 653
rect 451 643 453 651
rect 471 648 473 725
rect 571 725 613 727
rect 540 715 542 718
rect 571 715 573 725
rect 581 715 583 718
rect 591 715 593 718
rect 601 715 603 718
rect 540 693 542 707
rect 571 696 573 707
rect 581 692 583 707
rect 571 690 583 692
rect 540 686 542 689
rect 540 665 542 668
rect 461 646 473 648
rect 461 643 463 646
rect 540 643 542 657
rect 571 643 573 690
rect 591 687 593 707
rect 581 685 593 687
rect 581 643 583 685
rect 601 653 603 707
rect 591 651 603 653
rect 591 643 593 651
rect 611 648 613 725
rect 601 646 613 648
rect 601 643 603 646
rect 120 636 122 639
rect 151 623 153 639
rect 161 636 163 639
rect 171 615 173 639
rect 181 636 183 639
rect 260 636 262 639
rect 291 623 293 639
rect 301 636 303 639
rect 311 615 313 639
rect 321 636 323 639
rect 400 636 402 639
rect 431 623 433 639
rect 441 636 443 639
rect 451 615 453 639
rect 461 636 463 639
rect 540 636 542 639
rect 571 623 573 639
rect 581 636 583 639
rect 591 615 593 639
rect 601 636 603 639
<< polycontact >>
rect 27 1372 31 1376
rect 39 1365 43 1369
rect 57 1364 61 1368
rect 124 1372 128 1376
rect 155 1372 159 1376
rect 124 1322 128 1326
rect 165 1352 169 1356
rect 247 1372 251 1376
rect 259 1365 263 1369
rect 277 1364 281 1368
rect 344 1372 348 1376
rect 375 1372 379 1376
rect 344 1322 348 1326
rect 385 1352 389 1356
rect 467 1372 471 1376
rect 479 1365 483 1369
rect 497 1364 501 1368
rect 564 1372 568 1376
rect 595 1372 599 1376
rect 564 1322 568 1326
rect 605 1352 609 1356
rect 687 1372 691 1376
rect 699 1365 703 1369
rect 717 1364 721 1368
rect 784 1372 788 1376
rect 815 1372 819 1376
rect 784 1322 788 1326
rect 825 1352 829 1356
rect 155 1299 159 1303
rect 175 1291 179 1295
rect 375 1299 379 1303
rect 395 1291 399 1295
rect 595 1299 599 1303
rect 615 1291 619 1295
rect 815 1299 819 1303
rect 835 1291 839 1295
rect 230 1110 234 1114
rect 242 1103 246 1107
rect 260 1102 264 1106
rect 340 1110 344 1114
rect 352 1103 356 1107
rect 370 1102 374 1106
rect 489 1110 493 1114
rect 501 1103 505 1107
rect 519 1102 523 1106
rect 679 1110 683 1114
rect 691 1103 695 1107
rect 709 1102 713 1106
rect 340 1047 344 1051
rect 352 1040 356 1044
rect 364 1033 368 1037
rect 382 1035 386 1039
rect 489 1047 493 1051
rect 501 1040 505 1044
rect 513 1033 517 1037
rect 531 1035 535 1039
rect 679 1047 683 1051
rect 691 1040 695 1044
rect 703 1033 707 1037
rect 721 1035 725 1039
rect 489 977 493 981
rect 501 970 505 974
rect 513 963 517 967
rect 525 956 529 960
rect 543 962 547 966
rect 679 977 683 981
rect 691 970 695 974
rect 703 963 707 967
rect 715 956 719 960
rect 733 962 737 966
rect 679 900 683 904
rect 691 893 695 897
rect 703 886 707 890
rect 715 879 719 883
rect 727 872 731 876
rect 745 881 749 885
rect 231 808 235 812
rect 249 809 253 813
rect 261 816 265 820
rect 341 804 345 808
rect 359 802 363 806
rect 371 809 375 813
rect 383 816 387 820
rect 490 801 494 805
rect 508 795 512 799
rect 520 802 524 806
rect 532 809 536 813
rect 544 816 548 820
rect 680 797 684 801
rect 698 788 702 792
rect 710 795 714 799
rect 722 802 726 806
rect 734 809 738 813
rect 746 816 750 820
rect 116 696 120 700
rect 147 696 151 700
rect 116 646 120 650
rect 157 676 161 680
rect 256 696 260 700
rect 287 696 291 700
rect 256 646 260 650
rect 297 676 301 680
rect 396 696 400 700
rect 427 696 431 700
rect 396 646 400 650
rect 437 676 441 680
rect 536 696 540 700
rect 567 696 571 700
rect 536 646 540 650
rect 577 676 581 680
rect 147 623 151 627
rect 167 615 171 619
rect 287 623 291 627
rect 307 615 311 619
rect 427 623 431 627
rect 447 615 451 619
rect 567 623 571 627
rect 587 615 591 619
<< metal1 >>
rect -22 1148 -18 1429
rect -12 1397 895 1401
rect 24 1391 28 1397
rect 48 1391 52 1397
rect 56 1391 60 1397
rect 36 1376 40 1383
rect 15 1372 27 1376
rect 36 1372 52 1376
rect 6 1365 39 1369
rect 48 1368 52 1372
rect 64 1368 68 1383
rect 94 1372 98 1376
rect 48 1364 57 1368
rect 64 1364 72 1368
rect 48 1355 52 1364
rect 64 1355 68 1364
rect 108 1351 112 1397
rect 123 1391 127 1397
rect 153 1391 157 1397
rect 193 1391 197 1397
rect 244 1391 248 1397
rect 268 1391 272 1397
rect 276 1391 280 1397
rect 131 1376 135 1383
rect 120 1372 124 1376
rect 131 1372 155 1376
rect 131 1369 135 1372
rect 123 1361 127 1365
rect 117 1357 150 1361
rect 24 1311 28 1351
rect 56 1311 60 1351
rect 108 1347 141 1351
rect 123 1341 127 1347
rect 131 1326 135 1333
rect 86 1322 107 1326
rect 112 1322 124 1326
rect 131 1322 138 1326
rect 131 1319 135 1322
rect 123 1311 127 1315
rect 146 1311 150 1357
rect 158 1352 165 1356
rect 173 1350 177 1383
rect 256 1376 260 1383
rect 235 1372 247 1376
rect 256 1372 272 1376
rect 226 1365 259 1369
rect 268 1368 272 1372
rect 284 1368 288 1383
rect 314 1372 318 1376
rect 268 1364 277 1368
rect 284 1364 292 1368
rect 268 1355 272 1364
rect 284 1355 288 1364
rect 328 1351 332 1397
rect 343 1391 347 1397
rect 373 1391 377 1397
rect 413 1391 417 1397
rect 464 1391 468 1397
rect 488 1391 492 1397
rect 496 1391 500 1397
rect 351 1376 355 1383
rect 340 1372 344 1376
rect 351 1372 375 1376
rect 351 1369 355 1372
rect 343 1361 347 1365
rect 337 1357 370 1361
rect 173 1346 205 1350
rect 173 1319 177 1346
rect 153 1311 157 1315
rect 193 1311 197 1315
rect 244 1311 248 1351
rect 276 1311 280 1351
rect 328 1347 361 1351
rect 343 1341 347 1347
rect 351 1326 355 1333
rect 306 1322 327 1326
rect 332 1322 344 1326
rect 351 1322 358 1326
rect 351 1319 355 1322
rect 343 1311 347 1315
rect 366 1311 370 1357
rect 378 1352 385 1356
rect 393 1350 397 1383
rect 476 1376 480 1383
rect 455 1372 467 1376
rect 476 1372 492 1376
rect 446 1365 479 1369
rect 488 1368 492 1372
rect 504 1368 508 1383
rect 534 1372 538 1376
rect 488 1364 497 1368
rect 504 1364 512 1368
rect 488 1355 492 1364
rect 504 1355 508 1364
rect 548 1351 552 1397
rect 563 1391 567 1397
rect 593 1391 597 1397
rect 633 1391 637 1397
rect 684 1391 688 1397
rect 708 1391 712 1397
rect 716 1391 720 1397
rect 571 1376 575 1383
rect 560 1372 564 1376
rect 571 1372 595 1376
rect 571 1369 575 1372
rect 563 1361 567 1365
rect 557 1357 590 1361
rect 393 1346 425 1350
rect 393 1319 397 1346
rect 373 1311 377 1315
rect 413 1311 417 1315
rect 464 1311 468 1351
rect 496 1311 500 1351
rect 548 1347 581 1351
rect 563 1341 567 1347
rect 571 1326 575 1333
rect 526 1322 547 1326
rect 552 1322 564 1326
rect 571 1322 578 1326
rect 571 1319 575 1322
rect 563 1311 567 1315
rect 586 1311 590 1357
rect 598 1352 605 1356
rect 613 1350 617 1383
rect 696 1376 700 1383
rect 675 1372 687 1376
rect 696 1372 712 1376
rect 666 1365 699 1369
rect 708 1368 712 1372
rect 724 1368 728 1383
rect 754 1372 758 1376
rect 708 1364 717 1368
rect 724 1364 732 1368
rect 708 1355 712 1364
rect 724 1355 728 1364
rect 768 1351 772 1397
rect 783 1391 787 1397
rect 813 1391 817 1397
rect 853 1391 857 1397
rect 791 1376 795 1383
rect 780 1372 784 1376
rect 791 1372 815 1376
rect 791 1369 795 1372
rect 783 1361 787 1365
rect 777 1357 810 1361
rect 613 1346 645 1350
rect 613 1319 617 1346
rect 593 1311 597 1315
rect 633 1311 637 1315
rect 684 1311 688 1351
rect 716 1311 720 1351
rect 768 1347 801 1351
rect 783 1341 787 1347
rect 791 1326 795 1333
rect 746 1322 767 1326
rect 772 1322 784 1326
rect 791 1322 798 1326
rect 791 1319 795 1322
rect 783 1311 787 1315
rect 806 1311 810 1357
rect 818 1352 825 1356
rect 833 1350 837 1383
rect 833 1346 865 1350
rect 833 1319 837 1346
rect 813 1311 817 1315
rect 853 1311 857 1315
rect -12 1307 886 1311
rect 113 1299 155 1303
rect 333 1299 375 1303
rect 553 1299 595 1303
rect 773 1299 815 1303
rect 144 1291 175 1295
rect 364 1291 395 1295
rect 584 1291 615 1295
rect 804 1291 835 1295
rect 141 1216 661 1220
rect 666 1216 815 1220
rect 132 1207 798 1211
rect 803 1207 815 1211
rect 123 1198 471 1202
rect 476 1198 643 1202
rect 648 1198 815 1202
rect 114 1189 587 1193
rect 592 1189 652 1193
rect 657 1189 815 1193
rect 105 1180 322 1184
rect 327 1180 453 1184
rect 458 1180 624 1184
rect 629 1180 815 1184
rect 96 1171 417 1175
rect 422 1171 462 1175
rect 467 1171 634 1175
rect 639 1171 815 1175
rect 87 1162 212 1166
rect 217 1162 304 1166
rect 309 1162 435 1166
rect 440 1162 605 1166
rect 610 1162 815 1166
rect 78 1153 286 1157
rect 291 1153 313 1157
rect 318 1153 444 1157
rect 449 1153 614 1157
rect 619 1153 815 1157
rect -22 1144 73 1148
rect 78 1144 203 1148
rect 208 1144 295 1148
rect 300 1144 426 1148
rect 431 1144 596 1148
rect 601 1144 815 1148
rect 157 1135 895 1139
rect 82 744 86 1134
rect 100 743 104 1134
rect 118 752 122 1134
rect 136 761 140 1134
rect 157 1076 161 1135
rect 227 1129 231 1135
rect 251 1129 255 1135
rect 259 1129 263 1135
rect 337 1129 341 1135
rect 361 1129 365 1135
rect 369 1129 373 1135
rect 486 1129 490 1135
rect 510 1129 514 1135
rect 518 1129 522 1135
rect 676 1129 680 1135
rect 700 1129 704 1135
rect 708 1129 712 1135
rect 239 1114 243 1121
rect 218 1110 230 1114
rect 239 1110 255 1114
rect 209 1103 242 1107
rect 251 1106 255 1110
rect 267 1106 271 1121
rect 349 1114 353 1121
rect 328 1110 340 1114
rect 349 1110 365 1114
rect 251 1102 260 1106
rect 267 1102 277 1106
rect 251 1093 255 1102
rect 267 1093 271 1102
rect 319 1103 352 1107
rect 361 1106 365 1110
rect 377 1106 381 1121
rect 498 1114 502 1121
rect 477 1110 489 1114
rect 498 1110 514 1114
rect 361 1102 370 1106
rect 377 1102 408 1106
rect 361 1093 365 1102
rect 377 1093 381 1102
rect 468 1103 501 1107
rect 510 1106 514 1110
rect 526 1106 530 1121
rect 688 1114 692 1121
rect 667 1110 679 1114
rect 688 1110 704 1114
rect 510 1102 519 1106
rect 526 1102 578 1106
rect 510 1093 514 1102
rect 526 1093 530 1102
rect 658 1103 691 1107
rect 700 1106 704 1110
rect 716 1106 720 1121
rect 700 1102 709 1106
rect 716 1102 789 1106
rect 700 1093 704 1102
rect 716 1093 720 1102
rect 227 1085 231 1089
rect 259 1085 263 1089
rect 337 1085 341 1089
rect 369 1085 373 1089
rect 486 1085 490 1089
rect 518 1085 522 1089
rect 676 1085 680 1089
rect 708 1085 712 1089
rect 221 1081 886 1085
rect 157 1072 738 1076
rect 157 1006 161 1072
rect 337 1066 341 1072
rect 361 1066 365 1072
rect 381 1066 385 1072
rect 486 1066 490 1072
rect 510 1066 514 1072
rect 530 1066 534 1072
rect 676 1066 680 1072
rect 700 1066 704 1072
rect 720 1066 724 1072
rect 349 1051 353 1058
rect 373 1051 377 1058
rect 328 1047 340 1051
rect 349 1047 377 1051
rect 310 1040 352 1044
rect 373 1039 377 1047
rect 389 1039 393 1058
rect 498 1051 502 1058
rect 522 1051 526 1058
rect 477 1047 489 1051
rect 498 1047 526 1051
rect 459 1040 501 1044
rect 522 1039 526 1047
rect 538 1039 542 1058
rect 688 1051 692 1058
rect 712 1051 716 1058
rect 667 1047 679 1051
rect 688 1047 716 1051
rect 649 1040 691 1044
rect 712 1039 716 1047
rect 728 1039 732 1058
rect 301 1033 364 1037
rect 373 1035 382 1039
rect 389 1035 399 1039
rect 373 1023 377 1035
rect 389 1023 393 1035
rect 450 1033 513 1037
rect 522 1035 531 1039
rect 538 1035 569 1039
rect 522 1023 526 1035
rect 538 1023 542 1035
rect 640 1033 703 1037
rect 712 1035 721 1039
rect 728 1035 780 1039
rect 712 1023 716 1035
rect 728 1023 732 1035
rect 337 1015 341 1019
rect 381 1015 385 1019
rect 486 1015 490 1019
rect 530 1015 534 1019
rect 676 1015 680 1019
rect 720 1015 724 1019
rect 811 1015 815 1081
rect 331 1011 815 1015
rect 157 1002 750 1006
rect 157 929 161 1002
rect 486 996 490 1002
rect 510 996 514 1002
rect 534 996 538 1002
rect 542 996 546 1002
rect 676 996 680 1002
rect 700 996 704 1002
rect 724 996 728 1002
rect 732 996 736 1002
rect 498 981 502 988
rect 522 981 526 988
rect 477 977 489 981
rect 498 977 538 981
rect 459 970 501 974
rect 441 963 513 967
rect 534 966 538 977
rect 550 966 554 988
rect 688 981 692 988
rect 712 981 716 988
rect 667 977 679 981
rect 688 977 728 981
rect 649 970 691 974
rect 534 962 543 966
rect 550 962 560 966
rect 432 956 525 960
rect 534 946 538 962
rect 550 946 554 962
rect 630 963 703 967
rect 724 966 728 977
rect 740 966 744 988
rect 724 962 733 966
rect 740 962 771 966
rect 620 956 715 960
rect 724 946 728 962
rect 740 946 744 962
rect 486 938 490 942
rect 542 938 546 942
rect 676 938 680 942
rect 732 938 736 942
rect 811 938 815 1011
rect 480 934 815 938
rect 157 925 762 929
rect 157 845 161 925
rect 676 919 680 925
rect 700 919 704 925
rect 724 919 728 925
rect 744 919 748 925
rect 688 904 692 911
rect 712 904 716 911
rect 736 904 740 911
rect 667 900 679 904
rect 688 900 740 904
rect 649 893 691 897
rect 630 886 703 890
rect 736 885 740 900
rect 752 885 756 911
rect 611 879 715 883
rect 736 881 745 885
rect 752 881 762 885
rect 602 872 727 876
rect 736 862 740 881
rect 752 862 756 881
rect 676 854 680 858
rect 744 854 748 858
rect 811 854 815 934
rect 670 850 815 854
rect 157 841 759 845
rect 232 835 236 841
rect 264 835 268 841
rect 342 835 346 841
rect 386 835 390 841
rect 491 835 495 841
rect 547 835 551 841
rect 681 835 685 841
rect 749 835 753 841
rect 224 812 228 827
rect 240 812 244 827
rect 265 816 277 820
rect 218 808 228 812
rect 235 808 244 812
rect 253 809 286 813
rect 334 808 338 827
rect 350 808 354 827
rect 387 816 399 820
rect 375 809 408 813
rect 224 799 228 808
rect 240 806 244 808
rect 240 802 256 806
rect 329 804 338 808
rect 345 804 354 808
rect 252 799 256 802
rect 232 770 236 795
rect 240 770 244 795
rect 264 770 268 795
rect 334 792 338 804
rect 350 799 354 804
rect 363 802 417 806
rect 483 805 487 827
rect 499 805 503 827
rect 548 816 560 820
rect 536 809 569 813
rect 477 801 487 805
rect 494 801 503 805
rect 524 802 578 806
rect 673 801 677 827
rect 689 801 693 827
rect 750 816 762 820
rect 738 809 771 813
rect 726 802 780 806
rect 350 795 378 799
rect 350 792 354 795
rect 374 792 378 795
rect 342 770 346 788
rect 362 770 366 788
rect 386 770 390 788
rect 483 785 487 801
rect 499 792 503 801
rect 512 795 587 799
rect 667 797 677 801
rect 684 797 693 801
rect 499 788 539 792
rect 511 785 515 788
rect 535 785 539 788
rect 491 770 495 781
rect 499 770 503 781
rect 523 770 527 781
rect 547 770 551 781
rect 673 778 677 797
rect 689 785 693 797
rect 714 795 789 799
rect 702 788 798 792
rect 689 781 741 785
rect 689 778 693 781
rect 713 778 717 781
rect 737 778 741 781
rect 681 770 685 774
rect 701 770 705 774
rect 725 770 729 774
rect 749 770 753 774
rect 811 770 815 850
rect 218 766 815 770
rect 136 757 505 761
rect 118 748 365 752
rect 361 744 365 748
rect 501 744 505 757
rect 100 739 221 743
rect 88 721 895 725
rect 86 696 90 700
rect 100 675 104 721
rect 115 715 119 721
rect 145 715 149 721
rect 185 715 189 721
rect 123 700 127 707
rect 112 696 116 700
rect 123 696 147 700
rect 123 693 127 696
rect 115 685 119 689
rect 109 681 142 685
rect 100 671 133 675
rect 115 665 119 671
rect 123 650 127 657
rect 78 646 99 650
rect 104 646 116 650
rect 123 646 130 650
rect 123 643 127 646
rect 115 635 119 639
rect 138 635 142 681
rect 150 676 157 680
rect 165 674 169 707
rect 226 696 230 700
rect 240 675 244 721
rect 255 715 259 721
rect 285 715 289 721
rect 325 715 329 721
rect 263 700 267 707
rect 252 696 256 700
rect 263 696 287 700
rect 263 693 267 696
rect 255 685 259 689
rect 249 681 282 685
rect 165 670 197 674
rect 165 643 169 670
rect 240 671 273 675
rect 255 665 259 671
rect 263 650 267 657
rect 218 646 239 650
rect 244 646 256 650
rect 263 646 270 650
rect 263 643 267 646
rect 145 635 149 639
rect 185 635 189 639
rect 255 635 259 639
rect 278 635 282 681
rect 290 676 297 680
rect 305 674 309 707
rect 366 696 370 700
rect 380 675 384 721
rect 395 715 399 721
rect 425 715 429 721
rect 465 715 469 721
rect 403 700 407 707
rect 392 696 396 700
rect 403 696 427 700
rect 403 693 407 696
rect 395 685 399 689
rect 389 681 422 685
rect 305 670 337 674
rect 305 643 309 670
rect 380 671 413 675
rect 395 665 399 671
rect 403 650 407 657
rect 358 646 379 650
rect 384 646 396 650
rect 403 646 410 650
rect 403 643 407 646
rect 285 635 289 639
rect 325 635 329 639
rect 395 635 399 639
rect 418 635 422 681
rect 430 676 437 680
rect 445 674 449 707
rect 506 696 510 700
rect 520 675 524 721
rect 535 715 539 721
rect 565 715 569 721
rect 605 715 609 721
rect 543 700 547 707
rect 532 696 536 700
rect 543 696 567 700
rect 543 693 547 696
rect 535 685 539 689
rect 529 681 562 685
rect 445 670 477 674
rect 445 643 449 670
rect 520 671 553 675
rect 535 665 539 671
rect 543 650 547 657
rect 498 646 519 650
rect 524 646 536 650
rect 543 646 550 650
rect 543 643 547 646
rect 425 635 429 639
rect 465 635 469 639
rect 535 635 539 639
rect 558 635 562 681
rect 570 676 577 680
rect 585 674 589 707
rect 585 670 617 674
rect 585 643 589 670
rect 565 635 569 639
rect 605 635 609 639
rect 88 631 886 635
rect 105 623 147 627
rect 245 623 287 627
rect 385 623 427 627
rect 525 623 567 627
rect 136 615 167 619
rect 276 615 307 619
rect 416 615 447 619
rect 556 615 587 619
<< m2contact >>
rect 10 1372 15 1377
rect 1 1365 6 1370
rect 89 1372 94 1377
rect 98 1371 103 1376
rect 72 1363 77 1368
rect 115 1371 120 1376
rect 81 1322 86 1327
rect 107 1321 112 1326
rect 138 1321 143 1326
rect 153 1351 158 1356
rect 230 1372 235 1377
rect 221 1365 226 1370
rect 309 1372 314 1377
rect 318 1371 323 1376
rect 292 1363 297 1368
rect 335 1371 340 1376
rect 205 1345 210 1350
rect 301 1322 306 1327
rect 327 1321 332 1326
rect 358 1321 363 1326
rect 373 1351 378 1356
rect 450 1372 455 1377
rect 441 1365 446 1370
rect 529 1372 534 1377
rect 538 1371 543 1376
rect 512 1363 517 1368
rect 555 1371 560 1376
rect 425 1345 430 1350
rect 521 1322 526 1327
rect 547 1321 552 1326
rect 578 1321 583 1326
rect 593 1351 598 1356
rect 670 1372 675 1377
rect 661 1365 666 1370
rect 749 1372 754 1377
rect 758 1371 763 1376
rect 732 1363 737 1368
rect 895 1396 900 1401
rect 775 1371 780 1376
rect 645 1345 650 1350
rect 741 1322 746 1327
rect 767 1321 772 1326
rect 798 1321 803 1326
rect 813 1351 818 1356
rect 865 1345 870 1350
rect 886 1306 891 1311
rect 108 1299 113 1304
rect 328 1299 333 1304
rect 548 1299 553 1304
rect 768 1299 773 1304
rect 139 1291 144 1296
rect 359 1291 364 1296
rect 579 1291 584 1296
rect 799 1291 804 1296
rect 136 1216 141 1221
rect 661 1215 666 1220
rect 127 1207 132 1212
rect 798 1206 803 1211
rect 118 1198 123 1203
rect 471 1197 476 1202
rect 643 1197 648 1202
rect 109 1189 114 1194
rect 587 1188 592 1193
rect 652 1188 657 1193
rect 100 1180 105 1185
rect 322 1179 327 1184
rect 453 1179 458 1184
rect 624 1179 629 1184
rect 91 1171 96 1176
rect 417 1170 422 1175
rect 462 1170 467 1175
rect 634 1170 639 1175
rect 82 1162 87 1167
rect 212 1161 217 1166
rect 304 1161 309 1166
rect 435 1161 440 1166
rect 605 1161 610 1166
rect 73 1153 78 1158
rect 286 1152 291 1157
rect 313 1152 318 1157
rect 444 1152 449 1157
rect 614 1152 619 1157
rect 73 1143 78 1148
rect 203 1143 208 1148
rect 295 1144 300 1149
rect 426 1143 431 1148
rect 596 1143 601 1148
rect 82 1134 87 1139
rect 100 1134 105 1139
rect 118 1134 123 1139
rect 136 1134 141 1139
rect 81 739 86 744
rect 895 1134 900 1139
rect 213 1110 218 1115
rect 204 1103 209 1108
rect 323 1110 328 1115
rect 277 1101 282 1106
rect 314 1103 319 1108
rect 472 1110 477 1115
rect 408 1101 413 1106
rect 463 1103 468 1108
rect 662 1110 667 1115
rect 578 1101 583 1106
rect 653 1103 658 1108
rect 789 1101 794 1106
rect 323 1047 328 1052
rect 305 1040 310 1045
rect 472 1047 477 1052
rect 454 1040 459 1045
rect 662 1047 667 1052
rect 644 1040 649 1045
rect 296 1033 301 1038
rect 399 1034 404 1039
rect 445 1033 450 1038
rect 569 1034 574 1039
rect 635 1033 640 1038
rect 780 1034 785 1039
rect 886 1080 891 1085
rect 472 977 477 982
rect 454 970 459 975
rect 436 963 441 968
rect 662 977 667 982
rect 644 970 649 975
rect 427 956 432 961
rect 560 961 565 966
rect 625 963 630 968
rect 615 956 620 961
rect 771 961 776 966
rect 662 900 667 905
rect 644 893 649 898
rect 625 886 630 891
rect 606 879 611 884
rect 597 872 602 877
rect 762 880 767 885
rect 277 816 282 821
rect 213 807 218 812
rect 286 809 291 814
rect 399 816 404 821
rect 408 809 413 814
rect 324 803 329 808
rect 417 802 422 807
rect 560 816 565 821
rect 569 809 574 814
rect 472 800 477 805
rect 578 802 583 807
rect 762 816 767 821
rect 771 809 776 814
rect 780 802 785 807
rect 587 795 592 800
rect 662 796 667 801
rect 789 795 794 800
rect 798 788 803 793
rect 221 739 226 744
rect 361 739 366 744
rect 501 739 506 744
rect 895 721 900 726
rect 81 696 86 701
rect 90 695 95 700
rect 107 695 112 700
rect 73 646 78 651
rect 99 645 104 650
rect 130 645 135 650
rect 145 675 150 680
rect 221 696 226 701
rect 230 695 235 700
rect 247 695 252 700
rect 197 669 202 674
rect 213 646 218 651
rect 239 645 244 650
rect 270 645 275 650
rect 285 675 290 680
rect 361 696 366 701
rect 370 695 375 700
rect 387 695 392 700
rect 337 669 342 674
rect 353 646 358 651
rect 379 645 384 650
rect 410 645 415 650
rect 425 675 430 680
rect 501 696 506 701
rect 510 695 515 700
rect 527 695 532 700
rect 477 669 482 674
rect 493 646 498 651
rect 519 645 524 650
rect 550 645 555 650
rect 565 675 570 680
rect 617 669 622 674
rect 886 631 891 636
rect 100 623 105 628
rect 240 623 245 628
rect 380 623 385 628
rect 520 623 525 628
rect 131 615 136 620
rect 271 615 276 620
rect 411 615 416 620
rect 551 615 556 620
<< metal2 >>
rect 1 1412 89 1416
rect 221 1412 309 1416
rect 441 1412 529 1416
rect 661 1412 749 1416
rect 1 1370 5 1412
rect 10 1404 80 1408
rect 10 1377 14 1404
rect 73 1158 77 1363
rect 81 1327 85 1403
rect 89 1377 93 1412
rect 103 1371 115 1375
rect 99 1356 103 1371
rect 221 1370 225 1412
rect 230 1404 300 1408
rect 230 1377 234 1404
rect 99 1352 153 1356
rect 108 1304 112 1321
rect 139 1296 143 1321
rect 206 1283 210 1345
rect 82 1279 210 1283
rect 82 1167 86 1279
rect 293 1274 297 1363
rect 301 1327 305 1403
rect 309 1377 313 1412
rect 323 1371 335 1375
rect 319 1356 323 1371
rect 441 1370 445 1412
rect 450 1404 520 1408
rect 450 1377 454 1404
rect 319 1352 373 1356
rect 328 1304 332 1321
rect 359 1296 363 1321
rect 91 1270 297 1274
rect 91 1176 95 1270
rect 426 1265 430 1345
rect 100 1261 430 1265
rect 100 1185 104 1261
rect 513 1256 517 1363
rect 521 1327 525 1403
rect 529 1377 533 1412
rect 543 1371 555 1375
rect 539 1356 543 1371
rect 661 1370 665 1412
rect 670 1404 740 1408
rect 670 1377 674 1404
rect 539 1352 593 1356
rect 548 1304 552 1321
rect 579 1296 583 1321
rect 109 1252 517 1256
rect 109 1194 113 1252
rect 646 1247 650 1345
rect 118 1243 650 1247
rect 118 1203 122 1243
rect 733 1238 737 1363
rect 741 1327 745 1403
rect 749 1377 753 1412
rect 763 1371 775 1375
rect 759 1356 763 1371
rect 759 1352 813 1356
rect 768 1304 772 1321
rect 799 1296 803 1321
rect 127 1234 737 1238
rect 127 1212 131 1234
rect 866 1229 870 1345
rect 887 1311 891 1429
rect 896 1401 900 1429
rect 136 1225 870 1229
rect 136 1221 140 1225
rect 73 651 77 1143
rect 82 1139 86 1162
rect 100 1139 104 1180
rect 118 1139 122 1198
rect 136 1139 140 1216
rect 204 1108 208 1143
rect 213 1115 217 1161
rect 278 821 282 1101
rect 287 814 291 1152
rect 296 1038 300 1144
rect 305 1045 309 1161
rect 314 1108 318 1152
rect 323 1115 327 1179
rect 323 1052 327 1110
rect 400 821 404 1034
rect 409 814 413 1101
rect 81 701 85 739
rect 95 695 107 699
rect 91 680 95 695
rect 91 676 145 680
rect 100 628 104 645
rect 131 620 135 645
rect 198 601 202 669
rect 213 651 217 807
rect 418 807 422 1170
rect 427 961 431 1143
rect 436 968 440 1161
rect 445 1038 449 1152
rect 454 1045 458 1179
rect 463 1108 467 1170
rect 472 1115 476 1197
rect 472 1052 476 1110
rect 454 975 458 1040
rect 472 982 476 1047
rect 561 821 565 961
rect 570 814 574 1034
rect 579 807 583 1101
rect 324 743 328 803
rect 588 800 592 1188
rect 597 877 601 1143
rect 606 884 610 1161
rect 615 961 619 1152
rect 625 968 629 1179
rect 635 1038 639 1170
rect 644 1045 648 1197
rect 653 1108 657 1188
rect 662 1115 666 1215
rect 662 1052 666 1110
rect 644 975 648 1040
rect 662 982 666 1047
rect 625 891 629 963
rect 644 898 648 970
rect 662 905 666 977
rect 763 821 767 880
rect 772 814 776 961
rect 781 807 785 1034
rect 324 739 357 743
rect 221 701 225 739
rect 235 695 247 699
rect 231 680 235 695
rect 231 676 285 680
rect 240 628 244 645
rect 271 620 275 645
rect 338 601 342 669
rect 353 651 357 739
rect 472 743 476 800
rect 790 800 794 1101
rect 472 739 497 743
rect 361 701 365 739
rect 375 695 387 699
rect 371 680 375 695
rect 371 676 425 680
rect 380 628 384 645
rect 411 620 415 645
rect 478 601 482 669
rect 493 651 497 739
rect 501 701 505 739
rect 515 695 527 699
rect 511 680 515 695
rect 511 676 565 680
rect 520 628 524 645
rect 551 620 555 645
rect 618 601 622 669
rect 662 601 666 796
rect 799 793 803 1206
rect 887 1085 891 1306
rect 896 1139 900 1396
rect 887 636 891 1080
rect 896 726 900 1134
<< m3contact >>
rect 89 1412 94 1417
rect 309 1412 314 1417
rect 529 1412 534 1417
rect 749 1412 754 1417
rect 80 1403 85 1408
rect 300 1403 305 1408
rect 520 1403 525 1408
rect 740 1403 745 1408
<< metal3 >>
rect 80 1408 84 1429
rect 89 1417 93 1429
rect 300 1408 304 1429
rect 309 1417 313 1429
rect 520 1408 524 1429
rect 529 1417 533 1429
rect 740 1408 744 1429
rect 749 1417 753 1429
<< labels >>
rlabel metal1 -22 1425 -18 1429 4 c0
rlabel metal3 80 1425 84 1429 5 a0
rlabel metal3 89 1425 93 1429 5 b0
rlabel metal3 300 1425 304 1429 5 a1
rlabel metal3 309 1425 313 1429 5 b1
rlabel metal3 520 1425 524 1429 5 a2
rlabel metal3 529 1425 533 1429 5 b2
rlabel metal3 740 1425 744 1429 5 a3
rlabel metal3 749 1425 753 1429 5 b3
rlabel metal2 198 601 202 605 1 s0
rlabel metal2 338 601 342 605 1 s1
rlabel metal2 478 601 482 605 1 s2
rlabel metal2 618 601 622 605 1 s3
rlabel metal2 662 601 666 605 1 c4
rlabel metal2 887 1425 891 1429 5 gnd
rlabel metal2 896 1425 900 1429 6 vdd
<< end >>
