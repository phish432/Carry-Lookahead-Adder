magic
tech scmos
timestamp 1638827040
<< nwell >>
rect 64 -29 120 -9
rect 174 -29 230 -9
rect 323 -29 379 -9
rect 513 -29 569 -9
rect 174 -92 242 -72
rect 323 -92 391 -72
rect 513 -92 581 -72
rect 323 -162 403 -142
rect 513 -162 593 -142
rect 513 -239 605 -219
rect 61 -323 117 -303
rect 171 -323 239 -303
rect 320 -323 400 -303
rect 510 -323 602 -303
<< ntransistor >>
rect 77 -55 79 -51
rect 89 -55 91 -51
rect 107 -55 109 -51
rect 187 -55 189 -51
rect 199 -55 201 -51
rect 217 -55 219 -51
rect 336 -55 338 -51
rect 348 -55 350 -51
rect 366 -55 368 -51
rect 526 -55 528 -51
rect 538 -55 540 -51
rect 556 -55 558 -51
rect 187 -125 189 -121
rect 199 -125 201 -121
rect 211 -125 213 -121
rect 229 -125 231 -121
rect 336 -125 338 -121
rect 348 -125 350 -121
rect 360 -125 362 -121
rect 378 -125 380 -121
rect 526 -125 528 -121
rect 538 -125 540 -121
rect 550 -125 552 -121
rect 568 -125 570 -121
rect 336 -202 338 -198
rect 348 -202 350 -198
rect 360 -202 362 -198
rect 372 -202 374 -198
rect 390 -202 392 -198
rect 526 -202 528 -198
rect 538 -202 540 -198
rect 550 -202 552 -198
rect 562 -202 564 -198
rect 580 -202 582 -198
rect 526 -286 528 -282
rect 538 -286 540 -282
rect 550 -286 552 -282
rect 562 -286 564 -282
rect 574 -286 576 -282
rect 592 -286 594 -282
rect 72 -349 74 -345
rect 90 -349 92 -345
rect 102 -349 104 -345
rect 182 -356 184 -352
rect 200 -356 202 -352
rect 212 -356 214 -352
rect 224 -356 226 -352
rect 331 -363 333 -359
rect 349 -363 351 -359
rect 361 -363 363 -359
rect 373 -363 375 -359
rect 385 -363 387 -359
rect 521 -370 523 -366
rect 539 -370 541 -366
rect 551 -370 553 -366
rect 563 -370 565 -366
rect 575 -370 577 -366
rect 587 -370 589 -366
<< ptransistor >>
rect 77 -23 79 -15
rect 89 -23 91 -15
rect 107 -23 109 -15
rect 187 -23 189 -15
rect 199 -23 201 -15
rect 217 -23 219 -15
rect 336 -23 338 -15
rect 348 -23 350 -15
rect 366 -23 368 -15
rect 526 -23 528 -15
rect 538 -23 540 -15
rect 556 -23 558 -15
rect 187 -86 189 -78
rect 199 -86 201 -78
rect 211 -86 213 -78
rect 229 -86 231 -78
rect 336 -86 338 -78
rect 348 -86 350 -78
rect 360 -86 362 -78
rect 378 -86 380 -78
rect 526 -86 528 -78
rect 538 -86 540 -78
rect 550 -86 552 -78
rect 568 -86 570 -78
rect 336 -156 338 -148
rect 348 -156 350 -148
rect 360 -156 362 -148
rect 372 -156 374 -148
rect 390 -156 392 -148
rect 526 -156 528 -148
rect 538 -156 540 -148
rect 550 -156 552 -148
rect 562 -156 564 -148
rect 580 -156 582 -148
rect 526 -233 528 -225
rect 538 -233 540 -225
rect 550 -233 552 -225
rect 562 -233 564 -225
rect 574 -233 576 -225
rect 592 -233 594 -225
rect 72 -317 74 -309
rect 90 -317 92 -309
rect 102 -317 104 -309
rect 182 -317 184 -309
rect 200 -317 202 -309
rect 212 -317 214 -309
rect 224 -317 226 -309
rect 331 -317 333 -309
rect 349 -317 351 -309
rect 361 -317 363 -309
rect 373 -317 375 -309
rect 385 -317 387 -309
rect 521 -317 523 -309
rect 539 -317 541 -309
rect 551 -317 553 -309
rect 563 -317 565 -309
rect 575 -317 577 -309
rect 587 -317 589 -309
<< ndiffusion >>
rect 74 -55 77 -51
rect 79 -55 89 -51
rect 91 -55 94 -51
rect 106 -55 107 -51
rect 109 -55 110 -51
rect 184 -55 187 -51
rect 189 -55 199 -51
rect 201 -55 204 -51
rect 216 -55 217 -51
rect 219 -55 220 -51
rect 333 -55 336 -51
rect 338 -55 348 -51
rect 350 -55 353 -51
rect 365 -55 366 -51
rect 368 -55 369 -51
rect 523 -55 526 -51
rect 528 -55 538 -51
rect 540 -55 543 -51
rect 555 -55 556 -51
rect 558 -55 559 -51
rect 184 -125 187 -121
rect 189 -125 199 -121
rect 201 -125 211 -121
rect 213 -125 216 -121
rect 228 -125 229 -121
rect 231 -125 232 -121
rect 333 -125 336 -121
rect 338 -125 348 -121
rect 350 -125 360 -121
rect 362 -125 365 -121
rect 377 -125 378 -121
rect 380 -125 381 -121
rect 523 -125 526 -121
rect 528 -125 538 -121
rect 540 -125 550 -121
rect 552 -125 555 -121
rect 567 -125 568 -121
rect 570 -125 571 -121
rect 333 -202 336 -198
rect 338 -202 348 -198
rect 350 -202 360 -198
rect 362 -202 372 -198
rect 374 -202 377 -198
rect 389 -202 390 -198
rect 392 -202 393 -198
rect 523 -202 526 -198
rect 528 -202 538 -198
rect 540 -202 550 -198
rect 552 -202 562 -198
rect 564 -202 567 -198
rect 579 -202 580 -198
rect 582 -202 583 -198
rect 523 -286 526 -282
rect 528 -286 538 -282
rect 540 -286 550 -282
rect 552 -286 562 -282
rect 564 -286 574 -282
rect 576 -286 579 -282
rect 591 -286 592 -282
rect 594 -286 595 -282
rect 71 -349 72 -345
rect 74 -349 75 -345
rect 87 -349 90 -345
rect 92 -349 95 -345
rect 99 -349 102 -345
rect 104 -349 107 -345
rect 181 -356 182 -352
rect 184 -356 185 -352
rect 197 -356 200 -352
rect 202 -356 205 -352
rect 209 -356 212 -352
rect 214 -356 217 -352
rect 221 -356 224 -352
rect 226 -356 229 -352
rect 330 -363 331 -359
rect 333 -363 334 -359
rect 346 -363 349 -359
rect 351 -363 354 -359
rect 358 -363 361 -359
rect 363 -363 366 -359
rect 370 -363 373 -359
rect 375 -363 378 -359
rect 382 -363 385 -359
rect 387 -363 390 -359
rect 520 -370 521 -366
rect 523 -370 524 -366
rect 536 -370 539 -366
rect 541 -370 544 -366
rect 548 -370 551 -366
rect 553 -370 556 -366
rect 560 -370 563 -366
rect 565 -370 568 -366
rect 572 -370 575 -366
rect 577 -370 580 -366
rect 584 -370 587 -366
rect 589 -370 592 -366
<< pdiffusion >>
rect 74 -23 77 -15
rect 79 -23 82 -15
rect 86 -23 89 -15
rect 91 -23 94 -15
rect 106 -23 107 -15
rect 109 -23 110 -15
rect 184 -23 187 -15
rect 189 -23 192 -15
rect 196 -23 199 -15
rect 201 -23 204 -15
rect 216 -23 217 -15
rect 219 -23 220 -15
rect 333 -23 336 -15
rect 338 -23 341 -15
rect 345 -23 348 -15
rect 350 -23 353 -15
rect 365 -23 366 -15
rect 368 -23 369 -15
rect 523 -23 526 -15
rect 528 -23 531 -15
rect 535 -23 538 -15
rect 540 -23 543 -15
rect 555 -23 556 -15
rect 558 -23 559 -15
rect 184 -86 187 -78
rect 189 -86 192 -78
rect 196 -86 199 -78
rect 201 -86 204 -78
rect 208 -86 211 -78
rect 213 -86 216 -78
rect 228 -86 229 -78
rect 231 -86 232 -78
rect 333 -86 336 -78
rect 338 -86 341 -78
rect 345 -86 348 -78
rect 350 -86 353 -78
rect 357 -86 360 -78
rect 362 -86 365 -78
rect 377 -86 378 -78
rect 380 -86 381 -78
rect 523 -86 526 -78
rect 528 -86 531 -78
rect 535 -86 538 -78
rect 540 -86 543 -78
rect 547 -86 550 -78
rect 552 -86 555 -78
rect 567 -86 568 -78
rect 570 -86 571 -78
rect 333 -156 336 -148
rect 338 -156 341 -148
rect 345 -156 348 -148
rect 350 -156 353 -148
rect 357 -156 360 -148
rect 362 -156 365 -148
rect 369 -156 372 -148
rect 374 -156 377 -148
rect 389 -156 390 -148
rect 392 -156 393 -148
rect 523 -156 526 -148
rect 528 -156 531 -148
rect 535 -156 538 -148
rect 540 -156 543 -148
rect 547 -156 550 -148
rect 552 -156 555 -148
rect 559 -156 562 -148
rect 564 -156 567 -148
rect 579 -156 580 -148
rect 582 -156 583 -148
rect 523 -233 526 -225
rect 528 -233 531 -225
rect 535 -233 538 -225
rect 540 -233 543 -225
rect 547 -233 550 -225
rect 552 -233 555 -225
rect 559 -233 562 -225
rect 564 -233 567 -225
rect 571 -233 574 -225
rect 576 -233 579 -225
rect 591 -233 592 -225
rect 594 -233 595 -225
rect 71 -317 72 -309
rect 74 -317 75 -309
rect 87 -317 90 -309
rect 92 -317 102 -309
rect 104 -317 107 -309
rect 181 -317 182 -309
rect 184 -317 185 -309
rect 197 -317 200 -309
rect 202 -317 212 -309
rect 214 -317 224 -309
rect 226 -317 229 -309
rect 330 -317 331 -309
rect 333 -317 334 -309
rect 346 -317 349 -309
rect 351 -317 361 -309
rect 363 -317 373 -309
rect 375 -317 385 -309
rect 387 -317 390 -309
rect 520 -317 521 -309
rect 523 -317 524 -309
rect 536 -317 539 -309
rect 541 -317 551 -309
rect 553 -317 563 -309
rect 565 -317 575 -309
rect 577 -317 587 -309
rect 589 -317 592 -309
<< ndcontact >>
rect 70 -55 74 -51
rect 94 -55 98 -51
rect 102 -55 106 -51
rect 110 -55 114 -51
rect 180 -55 184 -51
rect 204 -55 208 -51
rect 212 -55 216 -51
rect 220 -55 224 -51
rect 329 -55 333 -51
rect 353 -55 357 -51
rect 361 -55 365 -51
rect 369 -55 373 -51
rect 519 -55 523 -51
rect 543 -55 547 -51
rect 551 -55 555 -51
rect 559 -55 563 -51
rect 180 -125 184 -121
rect 216 -125 220 -121
rect 224 -125 228 -121
rect 232 -125 236 -121
rect 329 -125 333 -121
rect 365 -125 369 -121
rect 373 -125 377 -121
rect 381 -125 385 -121
rect 519 -125 523 -121
rect 555 -125 559 -121
rect 563 -125 567 -121
rect 571 -125 575 -121
rect 329 -202 333 -198
rect 377 -202 381 -198
rect 385 -202 389 -198
rect 393 -202 397 -198
rect 519 -202 523 -198
rect 567 -202 571 -198
rect 575 -202 579 -198
rect 583 -202 587 -198
rect 519 -286 523 -282
rect 579 -286 583 -282
rect 587 -286 591 -282
rect 595 -286 599 -282
rect 67 -349 71 -345
rect 75 -349 79 -345
rect 83 -349 87 -345
rect 95 -349 99 -345
rect 107 -349 111 -345
rect 177 -356 181 -352
rect 185 -356 189 -352
rect 193 -356 197 -352
rect 205 -356 209 -352
rect 217 -356 221 -352
rect 229 -356 233 -352
rect 326 -363 330 -359
rect 334 -363 338 -359
rect 342 -363 346 -359
rect 354 -363 358 -359
rect 366 -363 370 -359
rect 378 -363 382 -359
rect 390 -363 394 -359
rect 516 -370 520 -366
rect 524 -370 528 -366
rect 532 -370 536 -366
rect 544 -370 548 -366
rect 556 -370 560 -366
rect 568 -370 572 -366
rect 580 -370 584 -366
rect 592 -370 596 -366
<< pdcontact >>
rect 70 -23 74 -15
rect 82 -23 86 -15
rect 94 -23 98 -15
rect 102 -23 106 -15
rect 110 -23 114 -15
rect 180 -23 184 -15
rect 192 -23 196 -15
rect 204 -23 208 -15
rect 212 -23 216 -15
rect 220 -23 224 -15
rect 329 -23 333 -15
rect 341 -23 345 -15
rect 353 -23 357 -15
rect 361 -23 365 -15
rect 369 -23 373 -15
rect 519 -23 523 -15
rect 531 -23 535 -15
rect 543 -23 547 -15
rect 551 -23 555 -15
rect 559 -23 563 -15
rect 180 -86 184 -78
rect 192 -86 196 -78
rect 204 -86 208 -78
rect 216 -86 220 -78
rect 224 -86 228 -78
rect 232 -86 236 -78
rect 329 -86 333 -78
rect 341 -86 345 -78
rect 353 -86 357 -78
rect 365 -86 369 -78
rect 373 -86 377 -78
rect 381 -86 385 -78
rect 519 -86 523 -78
rect 531 -86 535 -78
rect 543 -86 547 -78
rect 555 -86 559 -78
rect 563 -86 567 -78
rect 571 -86 575 -78
rect 329 -156 333 -148
rect 341 -156 345 -148
rect 353 -156 357 -148
rect 365 -156 369 -148
rect 377 -156 381 -148
rect 385 -156 389 -148
rect 393 -156 397 -148
rect 519 -156 523 -148
rect 531 -156 535 -148
rect 543 -156 547 -148
rect 555 -156 559 -148
rect 567 -156 571 -148
rect 575 -156 579 -148
rect 583 -156 587 -148
rect 519 -233 523 -225
rect 531 -233 535 -225
rect 543 -233 547 -225
rect 555 -233 559 -225
rect 567 -233 571 -225
rect 579 -233 583 -225
rect 587 -233 591 -225
rect 595 -233 599 -225
rect 67 -317 71 -309
rect 75 -317 79 -309
rect 83 -317 87 -309
rect 107 -317 111 -309
rect 177 -317 181 -309
rect 185 -317 189 -309
rect 193 -317 197 -309
rect 229 -317 233 -309
rect 326 -317 330 -309
rect 334 -317 338 -309
rect 342 -317 346 -309
rect 390 -317 394 -309
rect 516 -317 520 -309
rect 524 -317 528 -309
rect 532 -317 536 -309
rect 592 -317 596 -309
<< polysilicon >>
rect 77 -15 79 -12
rect 89 -15 91 -12
rect 107 -15 109 -12
rect 187 -15 189 -12
rect 199 -15 201 -12
rect 217 -15 219 -12
rect 336 -15 338 -12
rect 348 -15 350 -12
rect 366 -15 368 -12
rect 526 -15 528 -12
rect 538 -15 540 -12
rect 556 -15 558 -12
rect 77 -51 79 -23
rect 89 -51 91 -23
rect 107 -51 109 -23
rect 187 -51 189 -23
rect 199 -51 201 -23
rect 217 -51 219 -23
rect 336 -51 338 -23
rect 348 -51 350 -23
rect 366 -51 368 -23
rect 526 -51 528 -23
rect 538 -51 540 -23
rect 556 -51 558 -23
rect 77 -58 79 -55
rect 89 -58 91 -55
rect 107 -58 109 -55
rect 187 -58 189 -55
rect 199 -58 201 -55
rect 217 -58 219 -55
rect 336 -58 338 -55
rect 348 -58 350 -55
rect 366 -58 368 -55
rect 526 -58 528 -55
rect 538 -58 540 -55
rect 556 -58 558 -55
rect 187 -78 189 -75
rect 199 -78 201 -75
rect 211 -78 213 -75
rect 229 -78 231 -75
rect 336 -78 338 -75
rect 348 -78 350 -75
rect 360 -78 362 -75
rect 378 -78 380 -75
rect 526 -78 528 -75
rect 538 -78 540 -75
rect 550 -78 552 -75
rect 568 -78 570 -75
rect 187 -121 189 -86
rect 199 -121 201 -86
rect 211 -121 213 -86
rect 229 -121 231 -86
rect 336 -121 338 -86
rect 348 -121 350 -86
rect 360 -121 362 -86
rect 378 -121 380 -86
rect 526 -121 528 -86
rect 538 -121 540 -86
rect 550 -121 552 -86
rect 568 -121 570 -86
rect 187 -128 189 -125
rect 199 -128 201 -125
rect 211 -128 213 -125
rect 229 -128 231 -125
rect 336 -128 338 -125
rect 348 -128 350 -125
rect 360 -128 362 -125
rect 378 -128 380 -125
rect 526 -128 528 -125
rect 538 -128 540 -125
rect 550 -128 552 -125
rect 568 -128 570 -125
rect 336 -148 338 -145
rect 348 -148 350 -145
rect 360 -148 362 -145
rect 372 -148 374 -145
rect 390 -148 392 -145
rect 526 -148 528 -145
rect 538 -148 540 -145
rect 550 -148 552 -145
rect 562 -148 564 -145
rect 580 -148 582 -145
rect 336 -198 338 -156
rect 348 -198 350 -156
rect 360 -198 362 -156
rect 372 -198 374 -156
rect 390 -198 392 -156
rect 526 -198 528 -156
rect 538 -198 540 -156
rect 550 -198 552 -156
rect 562 -198 564 -156
rect 580 -198 582 -156
rect 336 -205 338 -202
rect 348 -205 350 -202
rect 360 -205 362 -202
rect 372 -205 374 -202
rect 390 -205 392 -202
rect 526 -205 528 -202
rect 538 -205 540 -202
rect 550 -205 552 -202
rect 562 -205 564 -202
rect 580 -205 582 -202
rect 526 -225 528 -222
rect 538 -225 540 -222
rect 550 -225 552 -222
rect 562 -225 564 -222
rect 574 -225 576 -222
rect 592 -225 594 -222
rect 526 -282 528 -233
rect 538 -282 540 -233
rect 550 -282 552 -233
rect 562 -282 564 -233
rect 574 -282 576 -233
rect 592 -282 594 -233
rect 526 -289 528 -286
rect 538 -289 540 -286
rect 550 -289 552 -286
rect 562 -289 564 -286
rect 574 -289 576 -286
rect 592 -289 594 -286
rect 72 -309 74 -306
rect 90 -309 92 -306
rect 102 -309 104 -306
rect 182 -309 184 -306
rect 200 -309 202 -306
rect 212 -309 214 -306
rect 224 -309 226 -306
rect 331 -309 333 -306
rect 349 -309 351 -306
rect 361 -309 363 -306
rect 373 -309 375 -306
rect 385 -309 387 -306
rect 521 -309 523 -306
rect 539 -309 541 -306
rect 551 -309 553 -306
rect 563 -309 565 -306
rect 575 -309 577 -306
rect 587 -309 589 -306
rect 72 -345 74 -317
rect 90 -345 92 -317
rect 102 -345 104 -317
rect 72 -352 74 -349
rect 90 -352 92 -349
rect 102 -352 104 -349
rect 182 -352 184 -317
rect 200 -352 202 -317
rect 212 -352 214 -317
rect 224 -352 226 -317
rect 182 -359 184 -356
rect 200 -359 202 -356
rect 212 -359 214 -356
rect 224 -359 226 -356
rect 331 -359 333 -317
rect 349 -359 351 -317
rect 361 -359 363 -317
rect 373 -359 375 -317
rect 385 -359 387 -317
rect 331 -366 333 -363
rect 349 -366 351 -363
rect 361 -366 363 -363
rect 373 -366 375 -363
rect 385 -366 387 -363
rect 521 -366 523 -317
rect 539 -366 541 -317
rect 551 -366 553 -317
rect 563 -366 565 -317
rect 575 -366 577 -317
rect 587 -366 589 -317
rect 521 -373 523 -370
rect 539 -373 541 -370
rect 551 -373 553 -370
rect 563 -373 565 -370
rect 575 -373 577 -370
rect 587 -373 589 -370
<< polycontact >>
rect 73 -34 77 -30
rect 85 -41 89 -37
rect 103 -42 107 -38
rect 183 -34 187 -30
rect 195 -41 199 -37
rect 213 -42 217 -38
rect 332 -34 336 -30
rect 344 -41 348 -37
rect 362 -42 366 -38
rect 522 -34 526 -30
rect 534 -41 538 -37
rect 552 -42 556 -38
rect 183 -97 187 -93
rect 195 -104 199 -100
rect 207 -111 211 -107
rect 225 -109 229 -105
rect 332 -97 336 -93
rect 344 -104 348 -100
rect 356 -111 360 -107
rect 374 -109 378 -105
rect 522 -97 526 -93
rect 534 -104 538 -100
rect 546 -111 550 -107
rect 564 -109 568 -105
rect 332 -167 336 -163
rect 344 -174 348 -170
rect 356 -181 360 -177
rect 368 -188 372 -184
rect 386 -182 390 -178
rect 522 -167 526 -163
rect 534 -174 538 -170
rect 546 -181 550 -177
rect 558 -188 562 -184
rect 576 -182 580 -178
rect 522 -244 526 -240
rect 534 -251 538 -247
rect 546 -258 550 -254
rect 558 -265 562 -261
rect 570 -272 574 -268
rect 588 -263 592 -259
rect 74 -336 78 -332
rect 92 -335 96 -331
rect 104 -328 108 -324
rect 184 -340 188 -336
rect 202 -342 206 -338
rect 214 -335 218 -331
rect 226 -328 230 -324
rect 333 -343 337 -339
rect 351 -349 355 -345
rect 363 -342 367 -338
rect 375 -335 379 -331
rect 387 -328 391 -324
rect 523 -347 527 -343
rect 541 -356 545 -352
rect 553 -349 557 -345
rect 565 -342 569 -338
rect 577 -335 581 -331
rect 589 -328 593 -324
<< metal1 >>
rect 0 72 504 76
rect 509 72 658 76
rect 0 63 641 67
rect 646 63 658 67
rect 0 54 314 58
rect 319 54 486 58
rect 491 54 658 58
rect 0 45 430 49
rect 435 45 495 49
rect 500 45 658 49
rect 0 36 165 40
rect 170 36 296 40
rect 301 36 467 40
rect 472 36 658 40
rect 0 27 260 31
rect 265 27 305 31
rect 310 27 477 31
rect 482 27 658 31
rect 0 18 55 22
rect 60 18 147 22
rect 152 18 278 22
rect 283 18 448 22
rect 453 18 658 22
rect 0 9 129 13
rect 134 9 156 13
rect 161 9 287 13
rect 292 9 457 13
rect 462 9 658 13
rect 0 0 46 4
rect 51 0 138 4
rect 143 0 269 4
rect 274 0 439 4
rect 444 0 658 4
rect 0 -9 569 -5
rect 0 -68 4 -9
rect 70 -15 74 -9
rect 94 -15 98 -9
rect 102 -15 106 -9
rect 180 -15 184 -9
rect 204 -15 208 -9
rect 212 -15 216 -9
rect 329 -15 333 -9
rect 353 -15 357 -9
rect 361 -15 365 -9
rect 519 -15 523 -9
rect 543 -15 547 -9
rect 551 -15 555 -9
rect 82 -30 86 -23
rect 61 -34 73 -30
rect 82 -34 98 -30
rect 52 -41 85 -37
rect 94 -38 98 -34
rect 110 -38 114 -23
rect 192 -30 196 -23
rect 171 -34 183 -30
rect 192 -34 208 -30
rect 94 -42 103 -38
rect 110 -42 120 -38
rect 94 -51 98 -42
rect 110 -51 114 -42
rect 162 -41 195 -37
rect 204 -38 208 -34
rect 220 -38 224 -23
rect 341 -30 345 -23
rect 320 -34 332 -30
rect 341 -34 357 -30
rect 204 -42 213 -38
rect 220 -42 251 -38
rect 204 -51 208 -42
rect 220 -51 224 -42
rect 311 -41 344 -37
rect 353 -38 357 -34
rect 369 -38 373 -23
rect 531 -30 535 -23
rect 510 -34 522 -30
rect 531 -34 547 -30
rect 353 -42 362 -38
rect 369 -42 421 -38
rect 353 -51 357 -42
rect 369 -51 373 -42
rect 501 -41 534 -37
rect 543 -38 547 -34
rect 559 -38 563 -23
rect 543 -42 552 -38
rect 559 -42 632 -38
rect 543 -51 547 -42
rect 559 -51 563 -42
rect 70 -59 74 -55
rect 102 -59 106 -55
rect 180 -59 184 -55
rect 212 -59 216 -55
rect 329 -59 333 -55
rect 361 -59 365 -55
rect 519 -59 523 -55
rect 551 -59 555 -55
rect 64 -63 658 -59
rect 0 -72 581 -68
rect 0 -138 4 -72
rect 180 -78 184 -72
rect 204 -78 208 -72
rect 224 -78 228 -72
rect 329 -78 333 -72
rect 353 -78 357 -72
rect 373 -78 377 -72
rect 519 -78 523 -72
rect 543 -78 547 -72
rect 563 -78 567 -72
rect 192 -93 196 -86
rect 216 -93 220 -86
rect 171 -97 183 -93
rect 192 -97 220 -93
rect 153 -104 195 -100
rect 216 -105 220 -97
rect 232 -105 236 -86
rect 341 -93 345 -86
rect 365 -93 369 -86
rect 320 -97 332 -93
rect 341 -97 369 -93
rect 302 -104 344 -100
rect 365 -105 369 -97
rect 381 -105 385 -86
rect 531 -93 535 -86
rect 555 -93 559 -86
rect 510 -97 522 -93
rect 531 -97 559 -93
rect 492 -104 534 -100
rect 555 -105 559 -97
rect 571 -105 575 -86
rect 144 -111 207 -107
rect 216 -109 225 -105
rect 232 -109 242 -105
rect 216 -121 220 -109
rect 232 -121 236 -109
rect 293 -111 356 -107
rect 365 -109 374 -105
rect 381 -109 412 -105
rect 365 -121 369 -109
rect 381 -121 385 -109
rect 483 -111 546 -107
rect 555 -109 564 -105
rect 571 -109 623 -105
rect 555 -121 559 -109
rect 571 -121 575 -109
rect 180 -129 184 -125
rect 224 -129 228 -125
rect 329 -129 333 -125
rect 373 -129 377 -125
rect 519 -129 523 -125
rect 563 -129 567 -125
rect 654 -129 658 -63
rect 174 -133 658 -129
rect 0 -142 593 -138
rect 0 -215 4 -142
rect 329 -148 333 -142
rect 353 -148 357 -142
rect 377 -148 381 -142
rect 385 -148 389 -142
rect 519 -148 523 -142
rect 543 -148 547 -142
rect 567 -148 571 -142
rect 575 -148 579 -142
rect 341 -163 345 -156
rect 365 -163 369 -156
rect 320 -167 332 -163
rect 341 -167 381 -163
rect 302 -174 344 -170
rect 284 -181 356 -177
rect 377 -178 381 -167
rect 393 -178 397 -156
rect 531 -163 535 -156
rect 555 -163 559 -156
rect 510 -167 522 -163
rect 531 -167 571 -163
rect 492 -174 534 -170
rect 377 -182 386 -178
rect 393 -182 403 -178
rect 275 -188 368 -184
rect 377 -198 381 -182
rect 393 -198 397 -182
rect 473 -181 546 -177
rect 567 -178 571 -167
rect 583 -178 587 -156
rect 567 -182 576 -178
rect 583 -182 614 -178
rect 463 -188 558 -184
rect 567 -198 571 -182
rect 583 -198 587 -182
rect 329 -206 333 -202
rect 385 -206 389 -202
rect 519 -206 523 -202
rect 575 -206 579 -202
rect 654 -206 658 -133
rect 323 -210 658 -206
rect 0 -219 605 -215
rect 0 -299 4 -219
rect 519 -225 523 -219
rect 543 -225 547 -219
rect 567 -225 571 -219
rect 587 -225 591 -219
rect 531 -240 535 -233
rect 555 -240 559 -233
rect 579 -240 583 -233
rect 510 -244 522 -240
rect 531 -244 583 -240
rect 492 -251 534 -247
rect 473 -258 546 -254
rect 579 -259 583 -244
rect 595 -259 599 -233
rect 454 -265 558 -261
rect 579 -263 588 -259
rect 595 -263 605 -259
rect 445 -272 570 -268
rect 579 -282 583 -263
rect 595 -282 599 -263
rect 519 -290 523 -286
rect 587 -290 591 -286
rect 654 -290 658 -210
rect 513 -294 658 -290
rect 0 -303 602 -299
rect 75 -309 79 -303
rect 107 -309 111 -303
rect 185 -309 189 -303
rect 229 -309 233 -303
rect 334 -309 338 -303
rect 390 -309 394 -303
rect 524 -309 528 -303
rect 592 -309 596 -303
rect 67 -332 71 -317
rect 83 -332 87 -317
rect 108 -328 120 -324
rect 61 -336 71 -332
rect 78 -336 87 -332
rect 96 -335 129 -331
rect 177 -336 181 -317
rect 193 -336 197 -317
rect 230 -328 242 -324
rect 218 -335 251 -331
rect 67 -345 71 -336
rect 83 -338 87 -336
rect 83 -342 99 -338
rect 172 -340 181 -336
rect 188 -340 197 -336
rect 95 -345 99 -342
rect 75 -374 79 -349
rect 83 -374 87 -349
rect 107 -374 111 -349
rect 177 -352 181 -340
rect 193 -345 197 -340
rect 206 -342 260 -338
rect 326 -339 330 -317
rect 342 -339 346 -317
rect 391 -328 403 -324
rect 379 -335 412 -331
rect 320 -343 330 -339
rect 337 -343 346 -339
rect 367 -342 421 -338
rect 516 -343 520 -317
rect 532 -343 536 -317
rect 593 -328 605 -324
rect 581 -335 614 -331
rect 569 -342 623 -338
rect 193 -349 221 -345
rect 193 -352 197 -349
rect 217 -352 221 -349
rect 185 -374 189 -356
rect 205 -374 209 -356
rect 229 -374 233 -356
rect 326 -359 330 -343
rect 342 -352 346 -343
rect 355 -349 430 -345
rect 510 -347 520 -343
rect 527 -347 536 -343
rect 342 -356 382 -352
rect 354 -359 358 -356
rect 378 -359 382 -356
rect 334 -374 338 -363
rect 342 -374 346 -363
rect 366 -374 370 -363
rect 390 -374 394 -363
rect 516 -366 520 -347
rect 532 -359 536 -347
rect 557 -349 632 -345
rect 545 -356 641 -352
rect 532 -363 584 -359
rect 532 -366 536 -363
rect 556 -366 560 -363
rect 580 -366 584 -363
rect 524 -374 528 -370
rect 544 -374 548 -370
rect 568 -374 572 -370
rect 592 -374 596 -370
rect 654 -374 658 -294
rect 61 -378 658 -374
<< m2contact >>
rect 504 71 509 76
rect 641 62 646 67
rect 314 53 319 58
rect 486 53 491 58
rect 430 44 435 49
rect 495 44 500 49
rect 165 35 170 40
rect 296 35 301 40
rect 467 35 472 40
rect 260 26 265 31
rect 305 26 310 31
rect 477 26 482 31
rect 55 17 60 22
rect 147 17 152 22
rect 278 17 283 22
rect 448 17 453 22
rect 129 8 134 13
rect 156 8 161 13
rect 287 8 292 13
rect 457 8 462 13
rect 46 -1 51 4
rect 138 0 143 5
rect 269 -1 274 4
rect 439 -1 444 4
rect 56 -34 61 -29
rect 47 -41 52 -36
rect 166 -34 171 -29
rect 120 -43 125 -38
rect 157 -41 162 -36
rect 315 -34 320 -29
rect 251 -43 256 -38
rect 306 -41 311 -36
rect 505 -34 510 -29
rect 421 -43 426 -38
rect 496 -41 501 -36
rect 632 -43 637 -38
rect 166 -97 171 -92
rect 148 -104 153 -99
rect 315 -97 320 -92
rect 297 -104 302 -99
rect 505 -97 510 -92
rect 487 -104 492 -99
rect 139 -111 144 -106
rect 242 -110 247 -105
rect 288 -111 293 -106
rect 412 -110 417 -105
rect 478 -111 483 -106
rect 623 -110 628 -105
rect 315 -167 320 -162
rect 297 -174 302 -169
rect 279 -181 284 -176
rect 505 -167 510 -162
rect 487 -174 492 -169
rect 270 -188 275 -183
rect 403 -183 408 -178
rect 468 -181 473 -176
rect 458 -188 463 -183
rect 614 -183 619 -178
rect 505 -244 510 -239
rect 487 -251 492 -246
rect 468 -258 473 -253
rect 449 -265 454 -260
rect 440 -272 445 -267
rect 605 -264 610 -259
rect 120 -328 125 -323
rect 56 -337 61 -332
rect 129 -335 134 -330
rect 242 -328 247 -323
rect 251 -335 256 -330
rect 167 -341 172 -336
rect 260 -342 265 -337
rect 403 -328 408 -323
rect 412 -335 417 -330
rect 315 -344 320 -339
rect 421 -342 426 -337
rect 605 -328 610 -323
rect 614 -335 619 -330
rect 623 -342 628 -337
rect 430 -349 435 -344
rect 505 -348 510 -343
rect 632 -349 637 -344
rect 641 -356 646 -351
<< metal2 >>
rect 47 -36 51 -1
rect 56 -29 60 17
rect 121 -323 125 -43
rect 130 -330 134 8
rect 139 -106 143 0
rect 148 -99 152 17
rect 157 -36 161 8
rect 166 -29 170 35
rect 166 -92 170 -34
rect 243 -323 247 -110
rect 252 -330 256 -43
rect 56 -390 60 -337
rect 261 -337 265 26
rect 270 -183 274 -1
rect 279 -176 283 17
rect 288 -106 292 8
rect 297 -99 301 35
rect 306 -36 310 26
rect 315 -29 319 53
rect 315 -92 319 -34
rect 297 -169 301 -104
rect 315 -162 319 -97
rect 404 -323 408 -183
rect 413 -330 417 -110
rect 422 -337 426 -43
rect 167 -390 171 -341
rect 431 -344 435 44
rect 440 -267 444 -1
rect 449 -260 453 17
rect 458 -183 462 8
rect 468 -176 472 35
rect 478 -106 482 26
rect 487 -99 491 53
rect 496 -36 500 44
rect 505 -29 509 71
rect 505 -92 509 -34
rect 487 -169 491 -104
rect 505 -162 509 -97
rect 468 -253 472 -181
rect 487 -246 491 -174
rect 505 -239 509 -167
rect 606 -323 610 -264
rect 615 -330 619 -183
rect 624 -337 628 -110
rect 315 -390 319 -344
rect 633 -344 637 -43
rect 505 -394 509 -348
rect 642 -351 646 62
<< labels >>
rlabel metal1 0 0 4 4 3 c0
rlabel metal1 0 9 4 13 3 g0
rlabel metal1 0 18 4 22 3 p0
rlabel metal1 0 27 4 31 3 g1
rlabel metal1 0 36 4 40 3 p1
rlabel metal1 0 45 4 49 3 g2
rlabel metal1 0 54 4 58 3 p2
rlabel metal1 0 63 4 67 3 g3
rlabel metal1 0 72 4 76 4 p3
rlabel metal2 56 -390 60 -386 1 c1
rlabel metal2 167 -390 171 -386 1 c2
rlabel metal2 315 -390 319 -386 1 c3
rlabel metal2 505 -394 509 -390 1 c4
rlabel metal1 61 -378 658 -374 1 gnd
rlabel metal1 0 -303 602 -299 1 vdd
rlabel metal1 0 -219 605 -215 1 vdd
rlabel metal1 0 -142 593 -138 1 vdd
rlabel metal1 0 -72 581 -68 1 vdd
rlabel metal1 0 -9 569 -5 1 vdd
rlabel metal1 64 -63 658 -59 1 gnd
rlabel metal1 174 -133 658 -129 1 gnd
rlabel metal1 323 -210 658 -206 1 gnd
rlabel metal1 513 -294 658 -290 1 gnd
<< end >>
