magic
tech scmos
timestamp 1638797210
<< nwell >>
rect 154 86 210 106
rect 253 86 277 106
rect 283 86 339 106
rect 374 86 430 106
rect 473 86 497 106
rect 503 86 559 106
rect 594 86 650 106
rect 693 86 717 106
rect 723 86 779 106
rect 814 86 870 106
rect 913 86 937 106
rect 943 86 999 106
rect 253 36 277 56
rect 473 36 497 56
rect 693 36 717 56
rect 913 36 937 56
<< ntransistor >>
rect 264 74 266 78
rect 167 60 169 64
rect 179 60 181 64
rect 197 60 199 64
rect 484 74 486 78
rect 387 60 389 64
rect 399 60 401 64
rect 417 60 419 64
rect 704 74 706 78
rect 607 60 609 64
rect 619 60 621 64
rect 637 60 639 64
rect 924 74 926 78
rect 827 60 829 64
rect 839 60 841 64
rect 857 60 859 64
rect 264 24 266 28
rect 295 24 297 28
rect 305 24 307 28
rect 315 24 317 28
rect 325 24 327 28
rect 484 24 486 28
rect 515 24 517 28
rect 525 24 527 28
rect 535 24 537 28
rect 545 24 547 28
rect 704 24 706 28
rect 735 24 737 28
rect 745 24 747 28
rect 755 24 757 28
rect 765 24 767 28
rect 924 24 926 28
rect 955 24 957 28
rect 965 24 967 28
rect 975 24 977 28
rect 985 24 987 28
<< ptransistor >>
rect 167 92 169 100
rect 179 92 181 100
rect 197 92 199 100
rect 264 92 266 100
rect 295 92 297 100
rect 305 92 307 100
rect 315 92 317 100
rect 325 92 327 100
rect 264 42 266 50
rect 387 92 389 100
rect 399 92 401 100
rect 417 92 419 100
rect 484 92 486 100
rect 515 92 517 100
rect 525 92 527 100
rect 535 92 537 100
rect 545 92 547 100
rect 484 42 486 50
rect 607 92 609 100
rect 619 92 621 100
rect 637 92 639 100
rect 704 92 706 100
rect 735 92 737 100
rect 745 92 747 100
rect 755 92 757 100
rect 765 92 767 100
rect 704 42 706 50
rect 827 92 829 100
rect 839 92 841 100
rect 857 92 859 100
rect 924 92 926 100
rect 955 92 957 100
rect 965 92 967 100
rect 975 92 977 100
rect 985 92 987 100
rect 924 42 926 50
<< ndiffusion >>
rect 263 74 264 78
rect 266 74 267 78
rect 164 60 167 64
rect 169 60 179 64
rect 181 60 184 64
rect 196 60 197 64
rect 199 60 200 64
rect 483 74 484 78
rect 486 74 487 78
rect 384 60 387 64
rect 389 60 399 64
rect 401 60 404 64
rect 416 60 417 64
rect 419 60 420 64
rect 703 74 704 78
rect 706 74 707 78
rect 604 60 607 64
rect 609 60 619 64
rect 621 60 624 64
rect 636 60 637 64
rect 639 60 640 64
rect 923 74 924 78
rect 926 74 927 78
rect 824 60 827 64
rect 829 60 839 64
rect 841 60 844 64
rect 856 60 857 64
rect 859 60 860 64
rect 263 24 264 28
rect 266 24 267 28
rect 293 24 295 28
rect 297 24 305 28
rect 307 24 309 28
rect 313 24 315 28
rect 317 24 325 28
rect 327 24 329 28
rect 483 24 484 28
rect 486 24 487 28
rect 513 24 515 28
rect 517 24 525 28
rect 527 24 529 28
rect 533 24 535 28
rect 537 24 545 28
rect 547 24 549 28
rect 703 24 704 28
rect 706 24 707 28
rect 733 24 735 28
rect 737 24 745 28
rect 747 24 749 28
rect 753 24 755 28
rect 757 24 765 28
rect 767 24 769 28
rect 923 24 924 28
rect 926 24 927 28
rect 953 24 955 28
rect 957 24 965 28
rect 967 24 969 28
rect 973 24 975 28
rect 977 24 985 28
rect 987 24 989 28
<< pdiffusion >>
rect 164 92 167 100
rect 169 92 172 100
rect 176 92 179 100
rect 181 92 184 100
rect 196 92 197 100
rect 199 92 200 100
rect 263 92 264 100
rect 266 92 267 100
rect 293 92 295 100
rect 297 92 305 100
rect 307 92 309 100
rect 313 92 315 100
rect 317 92 325 100
rect 327 92 329 100
rect 263 42 264 50
rect 266 42 267 50
rect 384 92 387 100
rect 389 92 392 100
rect 396 92 399 100
rect 401 92 404 100
rect 416 92 417 100
rect 419 92 420 100
rect 483 92 484 100
rect 486 92 487 100
rect 513 92 515 100
rect 517 92 525 100
rect 527 92 529 100
rect 533 92 535 100
rect 537 92 545 100
rect 547 92 549 100
rect 483 42 484 50
rect 486 42 487 50
rect 604 92 607 100
rect 609 92 612 100
rect 616 92 619 100
rect 621 92 624 100
rect 636 92 637 100
rect 639 92 640 100
rect 703 92 704 100
rect 706 92 707 100
rect 733 92 735 100
rect 737 92 745 100
rect 747 92 749 100
rect 753 92 755 100
rect 757 92 765 100
rect 767 92 769 100
rect 703 42 704 50
rect 706 42 707 50
rect 824 92 827 100
rect 829 92 832 100
rect 836 92 839 100
rect 841 92 844 100
rect 856 92 857 100
rect 859 92 860 100
rect 923 92 924 100
rect 926 92 927 100
rect 953 92 955 100
rect 957 92 965 100
rect 967 92 969 100
rect 973 92 975 100
rect 977 92 985 100
rect 987 92 989 100
rect 923 42 924 50
rect 926 42 927 50
<< ndcontact >>
rect 259 74 263 78
rect 267 74 271 78
rect 160 60 164 64
rect 184 60 188 64
rect 192 60 196 64
rect 200 60 204 64
rect 479 74 483 78
rect 487 74 491 78
rect 380 60 384 64
rect 404 60 408 64
rect 412 60 416 64
rect 420 60 424 64
rect 699 74 703 78
rect 707 74 711 78
rect 600 60 604 64
rect 624 60 628 64
rect 632 60 636 64
rect 640 60 644 64
rect 919 74 923 78
rect 927 74 931 78
rect 820 60 824 64
rect 844 60 848 64
rect 852 60 856 64
rect 860 60 864 64
rect 259 24 263 28
rect 267 24 271 28
rect 289 24 293 28
rect 309 24 313 28
rect 329 24 333 28
rect 479 24 483 28
rect 487 24 491 28
rect 509 24 513 28
rect 529 24 533 28
rect 549 24 553 28
rect 699 24 703 28
rect 707 24 711 28
rect 729 24 733 28
rect 749 24 753 28
rect 769 24 773 28
rect 919 24 923 28
rect 927 24 931 28
rect 949 24 953 28
rect 969 24 973 28
rect 989 24 993 28
<< pdcontact >>
rect 160 92 164 100
rect 172 92 176 100
rect 184 92 188 100
rect 192 92 196 100
rect 200 92 204 100
rect 259 92 263 100
rect 267 92 271 100
rect 289 92 293 100
rect 309 92 313 100
rect 329 92 333 100
rect 259 42 263 50
rect 267 42 271 50
rect 380 92 384 100
rect 392 92 396 100
rect 404 92 408 100
rect 412 92 416 100
rect 420 92 424 100
rect 479 92 483 100
rect 487 92 491 100
rect 509 92 513 100
rect 529 92 533 100
rect 549 92 553 100
rect 479 42 483 50
rect 487 42 491 50
rect 600 92 604 100
rect 612 92 616 100
rect 624 92 628 100
rect 632 92 636 100
rect 640 92 644 100
rect 699 92 703 100
rect 707 92 711 100
rect 729 92 733 100
rect 749 92 753 100
rect 769 92 773 100
rect 699 42 703 50
rect 707 42 711 50
rect 820 92 824 100
rect 832 92 836 100
rect 844 92 848 100
rect 852 92 856 100
rect 860 92 864 100
rect 919 92 923 100
rect 927 92 931 100
rect 949 92 953 100
rect 969 92 973 100
rect 989 92 993 100
rect 919 42 923 50
rect 927 42 931 50
<< polysilicon >>
rect 295 110 337 112
rect 167 100 169 103
rect 179 100 181 103
rect 197 100 199 103
rect 264 100 266 103
rect 295 100 297 110
rect 305 100 307 103
rect 315 100 317 103
rect 325 100 327 103
rect 167 64 169 92
rect 179 64 181 92
rect 197 64 199 92
rect 264 78 266 92
rect 295 81 297 92
rect 305 77 307 92
rect 295 75 307 77
rect 264 71 266 74
rect 167 57 169 60
rect 179 57 181 60
rect 197 57 199 60
rect 264 50 266 53
rect 264 28 266 42
rect 295 28 297 75
rect 315 72 317 92
rect 305 70 317 72
rect 305 28 307 70
rect 325 38 327 92
rect 315 36 327 38
rect 315 28 317 36
rect 335 33 337 110
rect 515 110 557 112
rect 387 100 389 103
rect 399 100 401 103
rect 417 100 419 103
rect 484 100 486 103
rect 515 100 517 110
rect 525 100 527 103
rect 535 100 537 103
rect 545 100 547 103
rect 387 64 389 92
rect 399 64 401 92
rect 417 64 419 92
rect 484 78 486 92
rect 515 81 517 92
rect 525 77 527 92
rect 515 75 527 77
rect 484 71 486 74
rect 387 57 389 60
rect 399 57 401 60
rect 417 57 419 60
rect 484 50 486 53
rect 325 31 337 33
rect 325 28 327 31
rect 484 28 486 42
rect 515 28 517 75
rect 535 72 537 92
rect 525 70 537 72
rect 525 28 527 70
rect 545 38 547 92
rect 535 36 547 38
rect 535 28 537 36
rect 555 33 557 110
rect 735 110 777 112
rect 607 100 609 103
rect 619 100 621 103
rect 637 100 639 103
rect 704 100 706 103
rect 735 100 737 110
rect 745 100 747 103
rect 755 100 757 103
rect 765 100 767 103
rect 607 64 609 92
rect 619 64 621 92
rect 637 64 639 92
rect 704 78 706 92
rect 735 81 737 92
rect 745 77 747 92
rect 735 75 747 77
rect 704 71 706 74
rect 607 57 609 60
rect 619 57 621 60
rect 637 57 639 60
rect 704 50 706 53
rect 545 31 557 33
rect 545 28 547 31
rect 704 28 706 42
rect 735 28 737 75
rect 755 72 757 92
rect 745 70 757 72
rect 745 28 747 70
rect 765 38 767 92
rect 755 36 767 38
rect 755 28 757 36
rect 775 33 777 110
rect 955 110 997 112
rect 827 100 829 103
rect 839 100 841 103
rect 857 100 859 103
rect 924 100 926 103
rect 955 100 957 110
rect 965 100 967 103
rect 975 100 977 103
rect 985 100 987 103
rect 827 64 829 92
rect 839 64 841 92
rect 857 64 859 92
rect 924 78 926 92
rect 955 81 957 92
rect 965 77 967 92
rect 955 75 967 77
rect 924 71 926 74
rect 827 57 829 60
rect 839 57 841 60
rect 857 57 859 60
rect 924 50 926 53
rect 765 31 777 33
rect 765 28 767 31
rect 924 28 926 42
rect 955 28 957 75
rect 975 72 977 92
rect 965 70 977 72
rect 965 28 967 70
rect 985 38 987 92
rect 975 36 987 38
rect 975 28 977 36
rect 995 33 997 110
rect 985 31 997 33
rect 985 28 987 31
rect 264 21 266 24
rect 295 8 297 24
rect 305 21 307 24
rect 315 0 317 24
rect 325 21 327 24
rect 484 21 486 24
rect 515 8 517 24
rect 525 21 527 24
rect 535 0 537 24
rect 545 21 547 24
rect 704 21 706 24
rect 735 8 737 24
rect 745 21 747 24
rect 755 0 757 24
rect 765 21 767 24
rect 924 21 926 24
rect 955 8 957 24
rect 965 21 967 24
rect 975 0 977 24
rect 985 21 987 24
<< polycontact >>
rect 163 81 167 85
rect 175 74 179 78
rect 193 73 197 77
rect 260 81 264 85
rect 291 81 295 85
rect 260 31 264 35
rect 301 61 305 65
rect 383 81 387 85
rect 395 74 399 78
rect 413 73 417 77
rect 480 81 484 85
rect 511 81 515 85
rect 480 31 484 35
rect 521 61 525 65
rect 603 81 607 85
rect 615 74 619 78
rect 633 73 637 77
rect 700 81 704 85
rect 731 81 735 85
rect 700 31 704 35
rect 741 61 745 65
rect 823 81 827 85
rect 835 74 839 78
rect 853 73 857 77
rect 920 81 924 85
rect 951 81 955 85
rect 920 31 924 35
rect 961 61 965 65
rect 291 8 295 12
rect 311 0 315 4
rect 511 8 515 12
rect 531 0 535 4
rect 731 8 735 12
rect 751 0 755 4
rect 951 8 955 12
rect 971 0 975 4
<< metal1 >>
rect 124 106 1031 110
rect 160 100 164 106
rect 184 100 188 106
rect 192 100 196 106
rect 172 85 176 92
rect 151 81 163 85
rect 172 81 188 85
rect 142 74 175 78
rect 184 77 188 81
rect 200 77 204 92
rect 230 81 234 85
rect 184 73 193 77
rect 200 73 208 77
rect 184 64 188 73
rect 200 64 204 73
rect 244 60 248 106
rect 259 100 263 106
rect 289 100 293 106
rect 329 100 333 106
rect 380 100 384 106
rect 404 100 408 106
rect 412 100 416 106
rect 267 85 271 92
rect 256 81 260 85
rect 267 81 291 85
rect 267 78 271 81
rect 259 70 263 74
rect 253 66 286 70
rect 160 20 164 60
rect 192 20 196 60
rect 244 56 277 60
rect 259 50 263 56
rect 267 35 271 42
rect 222 31 243 35
rect 248 31 260 35
rect 267 31 274 35
rect 267 28 271 31
rect 259 20 263 24
rect 282 20 286 66
rect 294 61 301 65
rect 309 59 313 92
rect 392 85 396 92
rect 371 81 383 85
rect 392 81 408 85
rect 362 74 395 78
rect 404 77 408 81
rect 420 77 424 92
rect 450 81 454 85
rect 404 73 413 77
rect 420 73 428 77
rect 404 64 408 73
rect 420 64 424 73
rect 464 60 468 106
rect 479 100 483 106
rect 509 100 513 106
rect 549 100 553 106
rect 600 100 604 106
rect 624 100 628 106
rect 632 100 636 106
rect 487 85 491 92
rect 476 81 480 85
rect 487 81 511 85
rect 487 78 491 81
rect 479 70 483 74
rect 473 66 506 70
rect 309 55 341 59
rect 309 28 313 55
rect 289 20 293 24
rect 329 20 333 24
rect 380 20 384 60
rect 412 20 416 60
rect 464 56 497 60
rect 479 50 483 56
rect 487 35 491 42
rect 442 31 463 35
rect 468 31 480 35
rect 487 31 494 35
rect 487 28 491 31
rect 479 20 483 24
rect 502 20 506 66
rect 514 61 521 65
rect 529 59 533 92
rect 612 85 616 92
rect 591 81 603 85
rect 612 81 628 85
rect 582 74 615 78
rect 624 77 628 81
rect 640 77 644 92
rect 670 81 674 85
rect 624 73 633 77
rect 640 73 648 77
rect 624 64 628 73
rect 640 64 644 73
rect 684 60 688 106
rect 699 100 703 106
rect 729 100 733 106
rect 769 100 773 106
rect 820 100 824 106
rect 844 100 848 106
rect 852 100 856 106
rect 707 85 711 92
rect 696 81 700 85
rect 707 81 731 85
rect 707 78 711 81
rect 699 70 703 74
rect 693 66 726 70
rect 529 55 561 59
rect 529 28 533 55
rect 509 20 513 24
rect 549 20 553 24
rect 600 20 604 60
rect 632 20 636 60
rect 684 56 717 60
rect 699 50 703 56
rect 707 35 711 42
rect 662 31 683 35
rect 688 31 700 35
rect 707 31 714 35
rect 707 28 711 31
rect 699 20 703 24
rect 722 20 726 66
rect 734 61 741 65
rect 749 59 753 92
rect 832 85 836 92
rect 811 81 823 85
rect 832 81 848 85
rect 802 74 835 78
rect 844 77 848 81
rect 860 77 864 92
rect 890 81 894 85
rect 844 73 853 77
rect 860 73 868 77
rect 844 64 848 73
rect 860 64 864 73
rect 904 60 908 106
rect 919 100 923 106
rect 949 100 953 106
rect 989 100 993 106
rect 927 85 931 92
rect 916 81 920 85
rect 927 81 951 85
rect 927 78 931 81
rect 919 70 923 74
rect 913 66 946 70
rect 749 55 781 59
rect 749 28 753 55
rect 729 20 733 24
rect 769 20 773 24
rect 820 20 824 60
rect 852 20 856 60
rect 904 56 937 60
rect 919 50 923 56
rect 927 35 931 42
rect 882 31 903 35
rect 908 31 920 35
rect 927 31 934 35
rect 927 28 931 31
rect 919 20 923 24
rect 942 20 946 66
rect 954 61 961 65
rect 969 59 973 92
rect 969 55 1001 59
rect 969 28 973 55
rect 949 20 953 24
rect 989 20 993 24
rect 124 16 1031 20
rect 249 8 291 12
rect 469 8 511 12
rect 689 8 731 12
rect 909 8 951 12
rect 280 0 311 4
rect 500 0 531 4
rect 720 0 751 4
rect 940 0 971 4
<< m2contact >>
rect 146 81 151 86
rect 137 74 142 79
rect 225 81 230 86
rect 234 80 239 85
rect 208 72 213 77
rect 251 80 256 85
rect 217 31 222 36
rect 243 30 248 35
rect 274 30 279 35
rect 289 60 294 65
rect 366 81 371 86
rect 357 74 362 79
rect 445 81 450 86
rect 454 80 459 85
rect 428 72 433 77
rect 471 80 476 85
rect 341 54 346 59
rect 437 31 442 36
rect 463 30 468 35
rect 494 30 499 35
rect 509 60 514 65
rect 586 81 591 86
rect 577 74 582 79
rect 665 81 670 86
rect 674 80 679 85
rect 648 72 653 77
rect 691 80 696 85
rect 561 54 566 59
rect 657 31 662 36
rect 683 30 688 35
rect 714 30 719 35
rect 729 60 734 65
rect 806 81 811 86
rect 797 74 802 79
rect 885 81 890 86
rect 894 80 899 85
rect 868 72 873 77
rect 911 80 916 85
rect 781 54 786 59
rect 877 31 882 36
rect 903 30 908 35
rect 934 30 939 35
rect 949 60 954 65
rect 1001 54 1006 59
rect 244 8 249 13
rect 464 8 469 13
rect 684 8 689 13
rect 904 8 909 13
rect 275 0 280 5
rect 495 0 500 5
rect 715 0 720 5
rect 935 0 940 5
<< metal2 >>
rect 137 121 225 125
rect 357 121 445 125
rect 577 121 665 125
rect 797 121 885 125
rect 137 79 141 121
rect 146 113 216 117
rect 146 86 150 113
rect 209 -12 213 72
rect 217 36 221 112
rect 225 86 229 121
rect 239 80 251 84
rect 235 65 239 80
rect 357 79 361 121
rect 366 113 436 117
rect 366 86 370 113
rect 235 61 289 65
rect 244 13 248 30
rect 275 5 279 30
rect 342 -12 346 54
rect 429 -12 433 72
rect 437 36 441 112
rect 445 86 449 121
rect 459 80 471 84
rect 455 65 459 80
rect 577 79 581 121
rect 586 113 656 117
rect 586 86 590 113
rect 455 61 509 65
rect 464 13 468 30
rect 495 5 499 30
rect 562 -12 566 54
rect 649 -12 653 72
rect 657 36 661 112
rect 665 86 669 121
rect 679 80 691 84
rect 675 65 679 80
rect 797 79 801 121
rect 806 113 876 117
rect 806 86 810 113
rect 675 61 729 65
rect 684 13 688 30
rect 715 5 719 30
rect 782 -12 786 54
rect 869 -12 873 72
rect 877 36 881 112
rect 885 86 889 121
rect 899 80 911 84
rect 895 65 899 80
rect 895 61 949 65
rect 904 13 908 30
rect 935 5 939 30
rect 1002 -12 1006 54
<< m3contact >>
rect 225 121 230 126
rect 445 121 450 126
rect 665 121 670 126
rect 885 121 890 126
rect 216 112 221 117
rect 436 112 441 117
rect 656 112 661 117
rect 876 112 881 117
<< metal3 >>
rect 216 117 220 138
rect 225 126 229 138
rect 436 117 440 138
rect 445 126 449 138
rect 656 117 660 138
rect 665 126 669 138
rect 876 117 880 138
rect 885 126 889 138
<< labels >>
rlabel metal3 216 134 220 138 5 a0
rlabel metal3 225 134 229 138 5 b0
rlabel metal3 436 134 440 138 5 a1
rlabel metal3 445 134 449 138 5 b1
rlabel metal3 656 134 660 138 5 a2
rlabel metal3 665 134 669 138 5 b2
rlabel metal3 876 134 880 138 5 a3
rlabel metal3 885 134 889 138 5 b3
rlabel metal1 124 106 1031 110 1 vdd
rlabel metal1 124 16 1031 20 1 gnd
rlabel metal2 209 -12 213 -8 1 g0
rlabel metal2 342 -12 346 -8 1 p0
rlabel metal2 429 -12 433 -8 1 g1
rlabel metal2 562 -12 566 -8 1 p1
rlabel metal2 649 -12 653 -8 1 g2
rlabel metal2 782 -12 786 -8 1 p2
rlabel metal2 869 -12 873 -8 1 g3
rlabel metal2 1002 -12 1006 -8 1 p3
<< end >>
