magic
tech scmos
timestamp 1638583042
<< nwell >>
rect 0 0 68 20
<< ntransistor >>
rect 13 -33 15 -29
rect 25 -33 27 -29
rect 37 -33 39 -29
rect 55 -33 57 -29
<< ptransistor >>
rect 13 6 15 14
rect 25 6 27 14
rect 37 6 39 14
rect 55 6 57 14
<< ndiffusion >>
rect 10 -33 13 -29
rect 15 -33 25 -29
rect 27 -33 37 -29
rect 39 -33 42 -29
rect 54 -33 55 -29
rect 57 -33 58 -29
<< pdiffusion >>
rect 10 6 13 14
rect 15 6 18 14
rect 22 6 25 14
rect 27 6 30 14
rect 34 6 37 14
rect 39 6 42 14
rect 54 6 55 14
rect 57 6 58 14
<< ndcontact >>
rect 6 -33 10 -29
rect 42 -33 46 -29
rect 50 -33 54 -29
rect 58 -33 62 -29
<< pdcontact >>
rect 6 6 10 14
rect 18 6 22 14
rect 30 6 34 14
rect 42 6 46 14
rect 50 6 54 14
rect 58 6 62 14
<< polysilicon >>
rect 13 14 15 17
rect 25 14 27 17
rect 37 14 39 17
rect 55 14 57 17
rect 13 -29 15 6
rect 25 -29 27 6
rect 37 -29 39 6
rect 55 -29 57 6
rect 13 -36 15 -33
rect 25 -36 27 -33
rect 37 -36 39 -33
rect 55 -36 57 -33
<< polycontact >>
rect 9 -5 13 -1
rect 21 -12 25 -8
rect 33 -19 37 -15
rect 51 -17 55 -13
<< metal1 >>
rect 0 20 68 24
rect 6 14 10 20
rect 30 14 34 20
rect 50 14 54 20
rect 18 -1 22 6
rect 42 -1 46 6
rect 0 -5 9 -1
rect 18 -5 46 -1
rect 0 -12 21 -8
rect 42 -13 46 -5
rect 58 -13 62 6
rect 0 -19 33 -15
rect 42 -17 51 -13
rect 58 -17 68 -13
rect 42 -29 46 -17
rect 58 -29 62 -17
rect 6 -37 10 -33
rect 50 -37 54 -33
rect 0 -41 68 -37
<< labels >>
rlabel metal1 0 -5 4 -1 3 in1
rlabel metal1 0 -12 4 -8 3 in2
rlabel metal1 0 -19 4 -15 3 in3
rlabel metal1 0 20 68 24 5 vdd
rlabel metal1 0 -41 68 -37 1 gnd
rlabel metal1 64 -17 68 -13 7 out
<< end >>
