* SPICE3 file created from or3.ext - technology: scmos

.option scale=0.09u

M1000 a_15_6# in1 vdd w_0_0# pfet w=8 l=2
+  ad=80 pd=36 as=96 ps=56
M1001 a_15_n33# in1 gnd Gnd nfet w=4 l=2
+  ad=68 pd=50 as=88 ps=68
M1002 a_27_6# in2 a_15_6# w_0_0# pfet w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1003 a_15_n33# in3 a_27_6# w_0_0# pfet w=8 l=2
+  ad=56 pd=30 as=0 ps=0
M1004 gnd in2 a_15_n33# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 out a_15_n33# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 a_15_n33# in3 gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 out a_15_n33# vdd w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
C0 out a_15_n33# 0.05fF
C1 a_15_n33# vdd 0.11fF
C2 w_0_0# out 0.03fF
C3 in1 in2 0.27fF
C4 w_0_0# vdd 0.12fF
C5 gnd out 0.08fF
C6 in1 vdd 0.02fF
C7 w_0_0# a_15_n33# 0.10fF
C8 in3 a_15_n33# 0.37fF
C9 gnd a_15_n33# 0.18fF
C10 in3 w_0_0# 0.06fF
C11 out vdd 0.11fF
C12 w_0_0# in1 0.06fF
C13 in3 in1 0.08fF
C14 a_15_n33# in2 0.08fF
C15 w_0_0# in2 0.06fF
C16 in3 in2 0.44fF
C17 gnd Gnd 0.28fF
C18 out Gnd 0.12fF
C19 vdd Gnd 0.16fF
C20 a_15_n33# Gnd 0.43fF
C21 in3 Gnd 0.34fF
C22 in2 Gnd 0.30fF
C23 in1 Gnd 0.27fF
C24 w_0_0# Gnd 1.37fF
