.include ../../TSMC_180nm.txt

** Parameters **
.param VSupply=1.8
.global vdd gnd

** Input Voltages **
VS vdd gnd VSupply

.param HIGH=VSupply
.param LOW=0

* A = a3 a2 a1 a0
VA0 a0 gnd pulse LOW  HIGH 0 100p 100p 40n 80n
VA1 a1 gnd pulse HIGH LOW  0 100p 100p 10n 20n
VA2 a2 gnd pulse HIGH LOW  0 100p 100p 20n 40n
VA3 a3 gnd pulse LOW  HIGH 0 100p 100p 20n 40n

* B = b3 b2 b1 b0
VB0 b0 gnd pulse HIGH LOW  0 100p 100p 40n 80n
VB1 b1 gnd pulse LOW  HIGH 0 100p 100p 20n 40n
VB2 b2 gnd pulse LOW  HIGH 0 100p 100p 10n 20n
VB3 b3 gnd pulse HIGH LOW  0 100p 100p 10n 20n

* Carry-In = c0
VC0 c0 gnd pulse HIGH LOW  0 100p 100p 20n 40n

** Circuit Description **
.option scale=0.09u

M1000 a_685_911# c0 vdd w_670_905# CMOSP w=8 l=2
+  ad=216 pd=102 as=4256 ps=2424
M1001 a_253_1351# a1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=1784 ps=1484
M1002 gnd a_339_785# a_334_788# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1003 a_33_1351# a0 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1004 a_381_1315# a1 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1005 a_685_1089# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1006 a_821_1315# a3 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1007 a_593_639# a_542_639# s3 Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1008 a_122_639# c0 vdd w_109_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1009 vdd a_116_696# a_346_1058# w_331_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=136 ps=66
M1010 vdd a_256_696# a_495_988# w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=160 ps=72
M1011 a_685_988# a_256_696# vdd w_670_982# CMOSP w=8 l=2
+  ad=160 pd=72 as=0 ps=0
M1012 a_698_827# a_696_771# a_678_771# w_667_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=56 ps=30
M1013 a_350_1315# a1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1014 a_570_1315# a2 vdd w_557_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1015 a_229_792# a_63_1351# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1016 a_503_1351# a_473_1383# vdd w_458_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1017 a_433_639# a_334_788# gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1018 vdd a_63_1351# a_346_1121# w_331_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1019 s0 c0 a_153_707# w_139_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1020 vdd a_396_696# a_685_1058# w_670_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=136 ps=66
M1021 a_313_707# a_256_696# s1 w_279_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1022 a_262_689# a_256_696# vdd w_249_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1023 a_339_785# a_369_785# gnd Gnd CMOSN w=4 l=2
+  ad=68 pd=50 as=0 ps=0
M1024 vdd a_130_1315# a_181_1383# w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1025 vdd a_570_1315# a_621_1383# w_587_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1026 a_495_988# a_396_696# vdd w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 vdd a_396_696# a_685_988# w_670_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 a_495_1019# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1029 vdd a_678_771# c4 w_667_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1030 a_253_1383# a1 vdd w_238_1377# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1031 vdd a_503_1351# a_685_1121# w_670_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1032 a_346_1121# a_63_1351# a_346_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=40 ps=28
M1033 a_346_1019# a_256_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1034 a_732_771# a_685_988# vdd w_670_982# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1035 a_253_1383# b1 a_253_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1036 a_693_1383# b3 a_693_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=40 ps=28
M1037 gnd a_542_778# a_488_778# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=80 ps=56
M1038 gnd a_229_792# a_224_795# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1039 a_381_1383# a_350_1365# vdd w_367_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1040 a_33_1383# a0 vdd w_18_1377# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1041 a_821_1383# a_790_1365# vdd w_807_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1042 gnd a_720_771# a_678_771# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=108 ps=78
M1043 a_520_827# a_518_778# a_508_827# w_477_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=80 ps=36
M1044 gnd a_402_689# a_453_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1045 a_130_1365# b0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1046 a_33_1383# b0 a_33_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1047 a_790_1365# b3 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1048 a_350_1365# b1 vdd w_337_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1049 a_685_1121# a_503_1351# a_685_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1050 a_685_1019# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1051 a_369_785# a_346_1121# vdd w_331_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1052 a_685_858# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1053 a_346_1058# c0 vdd w_331_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 a_153_639# c0 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1055 a_181_1315# a_130_1315# a_116_696# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1056 a_621_1315# a_570_1315# a_396_696# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1057 s1 a_256_696# a_293_639# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1058 a_593_707# a_536_696# s3 w_559_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1059 a_685_911# a_536_696# vdd w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 a_495_988# a_116_696# vdd w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 vdd a_63_1351# a_685_988# w_670_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 a_402_639# a_334_788# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1063 a_369_785# a_346_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1064 a_542_689# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1065 a_433_707# a_402_689# vdd w_419_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1066 gnd a_259_792# a_229_792# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 a_249_827# a_63_1351# a_229_792# w_218_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=56 ps=30
M1068 a_283_1351# a_253_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1069 a_236_1121# a_116_696# vdd w_221_1115# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1070 a_696_771# a_693_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1071 vdd b1 a_253_1383# w_238_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 vdd b3 a_693_1383# w_678_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1073 a_358_1019# a_116_696# a_346_1019# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1074 a_63_1351# a_33_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1075 gnd a_790_1365# a_841_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1076 a_236_1089# a_116_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1077 gnd a_122_689# a_173_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1078 a_381_785# a_346_1058# vdd w_331_1052# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1079 a_685_942# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1080 vdd a_488_778# a_483_781# w_477_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1081 vdd b0 a_33_1383# w_18_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 a_473_1351# a2 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1083 a_488_778# a_503_1351# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 a_709_858# a_256_696# a_697_858# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=40 ps=28
M1085 a_542_778# a_495_988# vdd w_480_982# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1086 s3 a_536_696# a_573_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1087 vdd a_229_792# a_224_795# w_218_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1088 a_181_1383# b0 a_116_696# w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1089 a_621_1383# b2 a_396_696# w_587_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1090 a_697_1019# a_396_696# a_685_1019# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1091 vdd a_381_785# a_371_827# w_328_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1092 a_122_639# c0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1093 a_678_771# a_732_771# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 a_685_911# a_256_696# vdd w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 a_601_1315# a2 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1096 vdd a_402_639# a_453_707# w_419_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1097 vdd a_256_696# a_495_1058# w_480_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=136 ps=66
M1098 a_262_689# a_256_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1099 a_153_707# a_122_689# vdd w_139_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 a_697_858# a_396_696# a_685_858# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 a_570_1315# a2 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1102 s1 a_224_795# a_293_707# w_279_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1103 a_130_1315# a0 vdd w_117_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1104 a_283_1351# a_253_1383# vdd w_238_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1105 a_790_1315# a3 vdd w_777_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1106 a_696_771# a_693_1383# vdd w_678_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1107 a_402_689# a_396_696# vdd w_389_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1108 vdd a_396_696# a_685_911# w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 vdd c0 a_236_1121# w_221_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 vdd a_283_1351# a_495_1121# w_480_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1111 vdd c0 a_495_988# w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 a_722_827# a_720_771# a_710_827# w_667_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=80 ps=36
M1113 a_63_1351# a_33_1383# vdd w_18_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1114 vdd a_790_1315# a_841_1383# w_807_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1115 a_507_942# a_256_696# a_495_942# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=40 ps=28
M1116 a_709_942# a_256_696# a_697_942# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=40 ps=28
M1117 vdd a_259_792# a_249_827# w_218_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 a_346_1058# c0 a_358_1019# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1119 a_116_696# b0 a_161_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1120 a_396_696# b2 a_601_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 a_473_1383# a2 vdd w_458_1377# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1122 a_236_1121# c0 a_236_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1123 a_495_1121# a_283_1351# a_495_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=40 ps=28
M1124 a_542_639# a_483_781# vdd w_529_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1125 a_453_639# a_402_639# s2 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1126 a_473_1383# b2 a_473_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1127 gnd a_542_689# a_593_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 vdd a_122_639# a_173_707# w_139_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1129 a_601_1383# a_570_1365# vdd w_587_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1130 a_495_942# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 a_697_942# a_396_696# a_685_942# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 gnd a_518_778# a_488_778# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 a_721_858# a_116_696# a_709_858# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1134 a_350_1365# b1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1135 s3 a_483_781# a_573_707# w_559_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1136 a_570_1365# b2 vdd w_557_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1137 a_259_792# a_236_1121# vdd w_221_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1138 a_518_778# a_495_1121# vdd w_480_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1139 a_495_1058# a_63_1351# vdd w_480_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 a_401_1315# a_350_1315# a_256_696# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1141 a_732_771# a_685_988# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1142 a_122_689# a_116_696# vdd w_109_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1143 gnd a_744_771# a_678_771# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 vdd a_116_696# a_685_911# w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 a_841_1315# a_790_1315# a_536_696# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1146 gnd a_381_785# a_339_785# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 a_381_785# a_346_1058# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1148 a_259_792# a_236_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1149 a_518_778# a_495_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1150 a_116_696# a0 a_161_1383# w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1151 a_396_696# a2 a_601_1383# w_587_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 a_708_771# a_685_1121# vdd w_670_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1153 a_685_1058# a_283_1351# vdd w_670_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 a_262_639# a_224_795# vdd w_249_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1155 a_173_639# a_122_639# s0 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1156 gnd a_262_689# a_313_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1157 a_532_827# a_530_778# a_520_827# w_477_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1158 vdd b2 a_473_1383# w_458_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 a_734_827# a_732_771# a_722_827# w_667_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1160 a_744_771# a_685_911# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1161 a_507_1019# a_256_696# a_495_1019# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1162 a_519_942# a_116_696# a_507_942# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1163 a_685_988# a_63_1351# a_709_942# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1164 a_708_771# a_685_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1165 a_573_639# a_483_781# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 gnd a_350_1365# a_401_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 a_744_771# a_685_911# vdd w_670_905# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1168 a_530_778# a_495_1058# vdd w_480_1052# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1169 a_693_1351# a3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 a_453_707# a_396_696# s2 w_419_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1171 gnd a_488_778# a_483_781# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1172 vdd a_542_639# a_593_707# w_559_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 a_401_1383# b1 a_256_696# w_367_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1174 a_841_1383# b3 a_536_696# w_807_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1175 a_402_689# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1176 a_161_1315# a0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 a_720_771# a_685_1058# vdd w_670_1052# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1178 a_678_771# a_708_771# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 a_359_827# a_283_1351# a_339_785# w_328_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=56 ps=30
M1180 a_790_1315# a3 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1181 a_130_1315# a0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1182 a_542_778# a_495_988# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1183 a_350_1315# a1 vdd w_337_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1184 a_293_639# a_224_795# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 vdd a_350_1315# a_401_1383# w_367_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 s2 a_396_696# a_433_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 gnd a_696_771# a_678_771# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 a_256_696# b1 a_381_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 a_495_1058# a_63_1351# a_507_1019# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1190 a_542_639# a_483_781# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1191 a_536_696# b3 a_821_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 a_173_707# a_116_696# s0 w_139_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 a_693_1383# a3 vdd w_678_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 vdd a_262_639# a_313_707# w_279_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 vdd a_339_785# a_334_788# w_328_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1196 vdd a_744_771# a_734_827# w_667_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 vdd a_542_778# a_532_827# w_477_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 a_495_988# c0 a_519_942# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1199 a_573_707# a_542_689# vdd w_559_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1200 a_122_689# a_116_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1201 a_161_1383# a_130_1365# vdd w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1202 a_570_1365# b2 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1203 a_685_1058# a_283_1351# a_697_1019# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1204 a_790_1365# b3 vdd w_777_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1205 a_130_1365# b0 vdd w_117_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1206 gnd a_678_771# c4 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1207 a_495_1058# a_396_696# vdd w_480_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 a_346_1058# a_256_696# vdd w_331_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 a_530_778# a_495_1058# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1210 s0 a_116_696# a_153_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 a_402_639# a_334_788# vdd w_389_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1212 a_371_827# a_369_785# a_359_827# w_328_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 gnd a_283_1351# a_339_785# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 a_256_696# a1 a_381_1383# w_367_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 a_495_1121# a_396_696# vdd w_480_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 a_685_988# a_536_696# vdd w_670_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 a_313_639# a_262_639# s1 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1218 a_262_639# a_224_795# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1219 a_536_696# a3 a_821_1383# w_807_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1220 a_346_1121# a_256_696# vdd w_331_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 a_503_1351# a_473_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1222 a_685_1058# a_536_696# vdd w_670_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 a_293_707# a_262_689# vdd w_279_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1224 a_720_771# a_685_1058# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1225 s2 a_334_788# a_433_707# w_419_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1226 a_495_1089# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 a_488_778# a_530_778# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 a_685_911# c0 a_721_858# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1229 gnd a_130_1365# a_181_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 gnd a_570_1365# a_621_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 a_346_1089# a_256_696# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 a_542_689# a_536_696# vdd w_529_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1233 a_685_1121# a_536_696# vdd w_670_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 a_710_827# a_708_771# a_698_827# w_667_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 a_508_827# a_503_1351# a_488_778# w_477_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=56 ps=30
C0 a_693_1383# w_678_1377# 0.09fF
C1 gnd a_402_689# 0.08fF
C2 a0 vdd 0.22fF
C3 a_283_1351# a_253_1383# 0.05fF
C4 a_283_1351# vdd 0.79fF
C5 a_495_1058# w_480_1052# 0.12fF
C6 a_536_696# a_685_988# 0.03fF
C7 a_262_639# vdd 0.11fF
C8 a_685_911# vdd 0.21fF
C9 gnd a_570_1315# 0.31fF
C10 a_536_696# c0 0.29fF
C11 gnd a_256_696# 0.85fF
C12 a_63_1351# w_670_982# 0.06fF
C13 a_536_696# a_396_696# 3.37fF
C14 a_503_1351# a_116_696# 0.17fF
C15 a_122_639# vdd 0.11fF
C16 a_530_778# a_503_1351# 0.08fF
C17 c0 w_109_651# 0.06fF
C18 a_122_639# a_122_689# 0.02fF
C19 a_542_689# vdd 0.74fF
C20 a_63_1351# vdd 1.05fF
C21 a_495_1121# w_480_1115# 0.09fF
C22 a_708_771# a_744_771# 0.08fF
C23 a_259_792# vdd 0.48fF
C24 gnd a0 0.76fF
C25 w_480_1052# a_256_696# 0.06fF
C26 a_283_1351# gnd 0.38fF
C27 w_670_982# a_732_771# 0.03fF
C28 a_503_1351# w_670_1115# 0.06fF
C29 w_117_1377# vdd 0.05fF
C30 a_346_1121# a_369_785# 0.05fF
C31 w_807_1377# a_790_1315# 0.06fF
C32 gnd a_262_639# 0.31fF
C33 vdd a_732_771# 0.11fF
C34 gnd a_685_911# 0.08fF
C35 a_283_1351# w_670_1052# 0.06fF
C36 b3 a_693_1383# 0.21fF
C37 b1 a_350_1365# 0.06fF
C38 a_495_1121# a_396_696# 0.03fF
C39 a_495_1058# a_396_696# 0.03fF
C40 a3 w_777_1327# 0.06fF
C41 s1 vdd 0.03fF
C42 w_419_701# a_396_696# 0.06fF
C43 a_224_795# a_256_696# 0.33fF
C44 a_116_696# w_139_701# 0.06fF
C45 a_693_1383# a3 0.03fF
C46 a_122_639# gnd 0.31fF
C47 a_346_1058# w_331_1052# 0.12fF
C48 a_570_1315# a2 0.36fF
C49 gnd a_542_689# 0.08fF
C50 a_63_1351# gnd 0.47fF
C51 a_402_689# a_396_696# 0.06fF
C52 gnd a_259_792# 0.17fF
C53 a_685_988# a_256_696# 0.08fF
C54 w_670_982# vdd 0.18fF
C55 w_328_821# a_283_1351# 0.06fF
C56 c0 a_256_696# 0.61fF
C57 a_518_778# vdd 0.45fF
C58 a_116_696# s0 0.12fF
C59 a_253_1383# vdd 0.05fF
C60 a_570_1315# a_396_696# 0.08fF
C61 a_495_988# vdd 0.10fF
C62 a_122_689# vdd 0.74fF
C63 w_587_1377# a_570_1315# 0.06fF
C64 a_63_1351# w_480_1052# 0.06fF
C65 gnd a_732_771# 0.25fF
C66 a_396_696# a_256_696# 3.67fF
C67 a_224_795# a_262_639# 0.36fF
C68 a_696_771# a_720_771# 0.08fF
C69 a_283_1351# w_480_1115# 0.06fF
C70 gnd s1 0.13fF
C71 b2 vdd 0.48fF
C72 a_685_1058# a_536_696# 0.03fF
C73 a_116_696# b0 0.12fF
C74 a_346_1121# w_331_1115# 0.09fF
C75 a_283_1351# c0 0.66fF
C76 a_283_1351# a_339_785# 0.37fF
C77 w_667_821# a_732_771# 0.06fF
C78 a_130_1365# a_130_1315# 0.02fF
C79 a_259_792# w_221_1115# 0.03fF
C80 c0 a_685_911# 0.11fF
C81 a_283_1351# a_396_696# 2.05fF
C82 gnd a_518_778# 0.34fF
C83 gnd a_253_1383# 0.04fF
C84 w_419_701# a_402_639# 0.06fF
C85 gnd vdd 14.37fF
C86 a_396_696# a_685_911# 0.17fF
C87 gnd a_495_988# 0.08fF
C88 a_63_1351# a_685_988# 0.11fF
C89 w_529_651# vdd 0.05fF
C90 a_122_639# c0 0.36fF
C91 a_122_689# gnd 0.08fF
C92 w_218_821# a_229_792# 0.10fF
C93 a_63_1351# c0 6.77fF
C94 a_536_696# a_503_1351# 0.83fF
C95 vdd w_670_1052# 0.14fF
C96 a_402_639# a_402_689# 0.02fF
C97 w_238_1377# a1 0.06fF
C98 b3 w_777_1377# 0.06fF
C99 b2 gnd 0.21fF
C100 w_667_821# vdd 0.15fF
C101 a_708_771# a_720_771# 1.45fF
C102 a_63_1351# a_396_696# 0.58fF
C103 w_480_1052# vdd 0.14fF
C104 w_117_1327# a0 0.06fF
C105 a_346_1058# a_116_696# 0.17fF
C106 a_685_988# a_732_771# 0.05fF
C107 a_542_778# w_477_821# 0.06fF
C108 w_279_701# a_256_696# 0.06fF
C109 a_488_778# w_477_821# 0.10fF
C110 a_116_696# a_130_1365# 0.08fF
C111 w_221_1115# vdd 0.14fF
C112 w_328_821# vdd 0.12fF
C113 a_708_771# a_685_1121# 0.05fF
C114 a_381_785# a_283_1351# 0.08fF
C115 a_224_795# vdd 0.22fF
C116 a_790_1315# vdd 0.11fF
C117 w_389_651# a_334_788# 0.06fF
C118 b3 a_790_1365# 0.06fF
C119 w_389_701# a_402_689# 0.03fF
C120 a_685_988# w_670_982# 0.11fF
C121 a_518_778# w_480_1115# 0.03fF
C122 w_480_1115# vdd 0.14fF
C123 a2 vdd 0.22fF
C124 a_685_988# vdd 0.10fF
C125 a_790_1365# a_536_696# 0.08fF
C126 s3 a_542_639# 0.08fF
C127 a_790_1365# a3 0.02fF
C128 a_339_785# vdd 0.11fF
C129 c0 vdd 6.36fF
C130 a_708_771# a_696_771# 1.90fF
C131 w_279_701# a_262_639# 0.06fF
C132 c0 a_495_988# 0.11fF
C133 a_396_696# w_670_982# 0.06fF
C134 a_122_689# c0 0.02fF
C135 a_283_1351# w_238_1377# 0.03fF
C136 a_685_1058# a_283_1351# 0.11fF
C137 b2 a2 0.97fF
C138 a_483_781# a_542_639# 0.36fF
C139 a_396_696# vdd 1.09fF
C140 a_396_696# a_495_988# 0.03fF
C141 a_503_1351# a_256_696# 6.82fF
C142 w_587_1377# vdd 0.11fF
C143 a_678_771# a_720_771# 0.08fF
C144 a_224_795# gnd 0.80fF
C145 gnd a_790_1315# 0.31fF
C146 a_542_778# w_480_982# 0.03fF
C147 w_249_701# a_262_689# 0.03fF
C148 b2 a_396_696# 0.12fF
C149 s3 w_559_701# 0.02fF
C150 b2 w_587_1377# 0.06fF
C151 a_530_778# w_477_821# 0.06fF
C152 a_685_1121# w_670_1115# 0.09fF
C153 a_116_696# w_670_905# 0.06fF
C154 a_116_696# w_331_1052# 0.06fF
C155 a_536_696# w_559_701# 0.06fF
C156 a_696_771# a_116_696# 0.09fF
C157 gnd a2 0.76fF
C158 gnd a_685_988# 0.08fF
C159 w_419_701# s2 0.02fF
C160 a_283_1351# a_503_1351# 0.17fF
C161 a_483_781# w_559_701# 0.06fF
C162 w_367_1377# a_350_1365# 0.19fF
C163 gnd a_339_785# 0.10fF
C164 gnd c0 1.30fF
C165 w_777_1327# vdd 0.05fF
C166 w_117_1327# vdd 0.05fF
C167 a_402_689# s2 0.08fF
C168 w_279_701# s1 0.02fF
C169 a_530_778# a_542_778# 0.69fF
C170 a_693_1383# vdd 0.05fF
C171 a_790_1365# w_807_1377# 0.19fF
C172 gnd a_396_696# 0.76fF
C173 a_350_1315# w_337_1327# 0.03fF
C174 a_236_1121# a_116_696# 0.03fF
C175 w_147_1377# b0 0.06fF
C176 b0 a_33_1383# 0.21fF
C177 a_530_778# a_488_778# 0.08fF
C178 vdd w_458_1377# 0.14fF
C179 a_116_696# a_130_1315# 0.08fF
C180 a_369_785# w_331_1115# 0.03fF
C181 a_396_696# w_670_1052# 0.06fF
C182 a_381_785# vdd 0.39fF
C183 a_350_1365# a1 0.02fF
C184 a_678_771# a_696_771# 0.70fF
C185 a_63_1351# a_503_1351# 0.17fF
C186 b2 w_458_1377# 0.06fF
C187 a_396_696# w_480_1052# 0.06fF
C188 w_279_701# vdd 0.11fF
C189 a_402_639# vdd 0.11fF
C190 w_678_1377# a_696_771# 0.03fF
C191 c0 w_221_1115# 0.06fF
C192 w_328_821# a_339_785# 0.10fF
C193 a_116_696# w_480_982# 0.06fF
C194 a_253_1383# w_238_1377# 0.09fF
C195 a_262_639# w_249_651# 0.03fF
C196 w_238_1377# vdd 0.14fF
C197 a_693_1383# gnd 0.04fF
C198 a_744_771# a_685_911# 0.05fF
C199 a_346_1121# a_256_696# 0.03fF
C200 a_685_1058# vdd 0.16fF
C201 w_337_1377# vdd 0.05fF
C202 a_224_795# a_396_696# 0.09fF
C203 a_256_696# a_350_1365# 0.08fF
C204 a_122_639# w_139_701# 0.06fF
C205 a_350_1315# w_367_1377# 0.06fF
C206 a_536_696# a_334_788# 0.09fF
C207 a_708_771# w_670_1115# 0.03fF
C208 a_381_785# gnd 0.17fF
C209 w_18_1377# b0 0.06fF
C210 a_396_696# w_480_1115# 0.06fF
C211 a_396_696# a_685_988# 0.17fF
C212 a_678_771# a_708_771# 0.08fF
C213 w_147_1377# a_130_1365# 0.19fF
C214 w_587_1377# a2 0.06fF
C215 b0 a0 0.97fF
C216 c0 a_396_696# 0.45fF
C217 w_389_701# vdd 0.05fF
C218 a_402_639# gnd 0.31fF
C219 a_518_778# a_503_1351# 1.59fF
C220 a_536_696# a_685_1121# 0.03fF
C221 a_122_639# s0 0.08fF
C222 a_350_1315# a1 0.36fF
C223 a_503_1351# vdd 0.62fF
C224 a_542_689# a_542_639# 0.02fF
C225 a_790_1315# w_777_1327# 0.03fF
C226 a_744_771# a_732_771# 0.52fF
C227 w_587_1377# a_396_696# 0.02fF
C228 a_685_1058# gnd 0.08fF
C229 w_419_701# a_334_788# 0.06fF
C230 w_777_1377# vdd 0.05fF
C231 a_346_1058# a_256_696# 0.03fF
C232 a_381_785# w_328_821# 0.06fF
C233 a_536_696# w_670_905# 0.06fF
C234 a_685_1058# w_670_1052# 0.12fF
C235 a_536_696# a_696_771# 7.08fF
C236 a_678_771# c4 0.05fF
C237 a_63_1351# a_346_1121# 0.21fF
C238 a3 a_696_771# 0.12fF
C239 a_483_781# w_477_821# 0.03fF
C240 a_402_689# a_334_788# 0.02fF
C241 a2 w_458_1377# 0.06fF
C242 a_542_689# w_559_701# 0.19fF
C243 a_350_1315# a_256_696# 0.08fF
C244 a_224_795# w_279_701# 0.06fF
C245 w_139_701# vdd 0.11fF
C246 gnd a_503_1351# 0.38fF
C247 w_249_651# vdd 0.05fF
C248 w_117_1377# b0 0.06fF
C249 a_262_689# a_256_696# 0.06fF
C250 a_122_689# w_139_701# 0.19fF
C251 a_744_771# vdd 0.13fF
C252 a_130_1365# a0 0.02fF
C253 a_488_778# a_483_781# 0.05fF
C254 a_790_1365# vdd 0.74fF
C255 vdd s2 0.03fF
C256 a_542_639# vdd 0.11fF
C257 b1 w_367_1377# 0.06fF
C258 s0 vdd 0.03fF
C259 a_122_689# s0 0.08fF
C260 a_262_689# a_262_639# 0.02fF
C261 a_346_1121# vdd 0.05fF
C262 w_147_1377# a_130_1315# 0.06fF
C263 b0 vdd 0.48fF
C264 b1 a1 0.97fF
C265 vdd a_350_1365# 0.74fF
C266 gnd a_744_771# 0.17fF
C267 a_685_1058# a_396_696# 0.17fF
C268 w_559_701# vdd 0.11fF
C269 w_670_905# a_256_696# 0.06fF
C270 w_331_1052# a_256_696# 0.06fF
C271 a_696_771# a_256_696# 0.09fF
C272 a_790_1365# gnd 0.08fF
C273 gnd s2 0.13fF
C274 w_117_1377# a_130_1365# 0.03fF
C275 a_503_1351# a2 0.12fF
C276 gnd a_542_639# 0.31fF
C277 a_744_771# w_667_821# 0.06fF
C278 gnd s0 0.13fF
C279 a_536_696# a_116_696# 0.25fF
C280 a_542_639# w_529_651# 0.03fF
C281 c0 a_503_1351# 0.75fF
C282 w_389_701# a_396_696# 0.06fF
C283 a_116_696# w_109_701# 0.06fF
C284 a_283_1351# a_696_771# 0.09fF
C285 a_503_1351# a_396_696# 7.17fF
C286 b1 a_256_696# 0.12fF
C287 a_720_771# a_732_771# 1.00fF
C288 a_63_1351# a_229_792# 0.21fF
C289 gnd a_346_1121# 0.08fF
C290 a_570_1365# w_557_1377# 0.03fF
C291 gnd b0 0.21fF
C292 a_536_696# w_670_1115# 0.06fF
C293 a_685_911# w_670_905# 0.14fF
C294 a_262_689# s1 0.08fF
C295 a_346_1058# vdd 0.16fF
C296 gnd a_350_1365# 0.08fF
C297 a_224_795# w_249_651# 0.06fF
C298 a_473_1383# vdd 0.05fF
C299 a_116_696# w_147_1377# 0.02fF
C300 a_790_1365# a_790_1315# 0.02fF
C301 a_530_778# a_495_1058# 0.05fF
C302 a_130_1365# vdd 0.74fF
C303 b3 w_678_1377# 0.06fF
C304 a0 a_130_1315# 0.36fF
C305 a_283_1351# a_369_785# 1.29fF
C306 a_350_1315# vdd 0.11fF
C307 a_63_1351# a_696_771# 0.09fF
C308 c0 w_139_701# 0.06fF
C309 b2 a_473_1383# 0.21fF
C310 a_256_696# w_480_982# 0.06fF
C311 a3 w_678_1377# 0.06fF
C312 a_720_771# vdd 0.11fF
C313 a_262_689# vdd 0.74fF
C314 vdd a_334_788# 0.22fF
C315 a_63_1351# w_218_821# 0.06fF
C316 a_503_1351# w_458_1377# 0.03fF
C317 a_696_771# a_732_771# 0.08fF
C318 a_346_1058# gnd 0.08fF
C319 w_218_821# a_259_792# 0.06fF
C320 a_259_792# a_236_1121# 0.05fF
C321 a_570_1315# w_557_1327# 0.03fF
C322 a_396_696# s2 0.12fF
C323 a_116_696# a_256_696# 2.73fF
C324 a_473_1383# gnd 0.04fF
C325 a_229_792# vdd 0.11fF
C326 w_331_1115# a_256_696# 0.06fF
C327 a_685_1121# vdd 0.05fF
C328 gnd a_130_1365# 0.08fF
C329 a_350_1315# gnd 0.31fF
C330 a_518_778# w_477_821# 0.06fF
C331 gnd a_262_689# 0.08fF
C332 gnd a_720_771# 0.34fF
C333 w_477_821# vdd 0.14fF
C334 a_283_1351# a_116_696# 6.72fF
C335 gnd a_334_788# 0.89fF
C336 w_670_905# vdd 0.19fF
C337 w_331_1052# vdd 0.14fF
C338 a_696_771# vdd 0.20fF
C339 a_720_771# w_670_1052# 0.03fF
C340 b3 a_536_696# 0.12fF
C341 b3 a3 0.97fF
C342 a_116_696# a_685_911# 0.08fF
C343 s3 a_536_696# 0.12fF
C344 a_720_771# w_667_821# 0.06fF
C345 w_249_701# a_256_696# 0.06fF
C346 a_570_1315# a_570_1365# 0.02fF
C347 a_518_778# a_542_778# 0.08fF
C348 a_708_771# a_732_771# 0.08fF
C349 gnd a_229_792# 0.05fF
C350 a_542_778# vdd 0.30fF
C351 w_337_1327# a1 0.06fF
C352 w_218_821# vdd 0.11fF
C353 a_542_778# a_495_988# 0.05fF
C354 a_488_778# a_518_778# 0.08fF
C355 gnd a_685_1121# 0.08fF
C356 a_488_778# vdd 0.11fF
C357 a_236_1121# vdd 0.05fF
C358 a_536_696# a_483_781# 0.32fF
C359 b1 a_253_1383# 0.21fF
C360 a_369_785# vdd 0.45fF
C361 a_63_1351# a_116_696# 7.59fF
C362 b1 vdd 0.48fF
C363 a_130_1315# vdd 0.11fF
C364 a_63_1351# w_331_1115# 0.06fF
C365 a_473_1383# a2 0.03fF
C366 a_346_1058# c0 0.11fF
C367 w_328_821# a_334_788# 0.03fF
C368 a_224_795# a_262_689# 0.02fF
C369 a_402_639# s2 0.08fF
C370 gnd a_696_771# 0.47fF
C371 a_708_771# vdd 0.11fF
C372 gnd a_542_778# 0.17fF
C373 vdd w_480_982# 0.18fF
C374 a_224_795# a_229_792# 0.05fF
C375 a_696_771# w_667_821# 0.06fF
C376 a_495_988# w_480_982# 0.11fF
C377 b3 w_807_1377# 0.06fF
C378 gnd a_488_778# 0.11fF
C379 a_339_785# a_334_788# 0.05fF
C380 w_367_1377# a1 0.06fF
C381 gnd a_236_1121# 0.08fF
C382 gnd a_369_785# 0.25fF
C383 gnd b1 0.21fF
C384 a_536_696# w_807_1377# 0.02fF
C385 gnd a_130_1315# 0.31fF
C386 a3 w_807_1377# 0.06fF
C387 a_396_696# a_334_788# 0.32fF
C388 w_389_651# vdd 0.05fF
C389 a_536_696# w_529_701# 0.06fF
C390 a_678_771# a_732_771# 0.08fF
C391 c4 vdd 0.20fF
C392 a_530_778# a_518_778# 1.15fF
C393 a_116_696# vdd 1.21fF
C394 a_530_778# vdd 0.37fF
C395 a_116_696# a_495_988# 0.08fF
C396 a_536_696# a_256_696# 0.41fF
C397 w_331_1115# vdd 0.14fF
C398 w_337_1377# a_350_1365# 0.03fF
C399 a_122_689# a_116_696# 0.06fF
C400 w_557_1327# vdd 0.05fF
C401 a_708_771# gnd 0.42fF
C402 a_473_1383# w_458_1377# 0.09fF
C403 a_790_1365# w_777_1377# 0.03fF
C404 a_381_785# a_346_1058# 0.05fF
C405 w_367_1377# a_256_696# 0.02fF
C406 w_419_701# a_402_689# 0.19fF
C407 a_236_1121# w_221_1115# 0.09fF
C408 a_224_795# w_218_821# 0.03fF
C409 w_670_1115# vdd 0.14fF
C410 w_328_821# a_369_785# 0.06fF
C411 c0 w_670_905# 0.06fF
C412 c0 w_331_1052# 0.06fF
C413 a_696_771# c0 0.09fF
C414 a_708_771# w_667_821# 0.06fF
C415 a_536_696# a_283_1351# 0.33fF
C416 a_678_771# vdd 0.11fF
C417 a_396_696# w_670_905# 0.06fF
C418 a_495_1058# a_256_696# 0.17fF
C419 a_696_771# a_396_696# 6.93fF
C420 a_536_696# a_685_911# 0.03fF
C421 w_249_701# vdd 0.05fF
C422 gnd c4 0.25fF
C423 gnd a_116_696# 0.85fF
C424 a_530_778# gnd 0.25fF
C425 w_678_1377# vdd 0.14fF
C426 c0 a_236_1121# 0.21fF
C427 a_570_1365# vdd 0.74fF
C428 w_139_701# s0 0.02fF
C429 w_18_1377# a_33_1383# 0.09fF
C430 a_339_785# a_369_785# 0.08fF
C431 s3 a_542_689# 0.08fF
C432 w_147_1377# a0 0.06fF
C433 w_279_701# a_262_689# 0.19fF
C434 a_33_1383# a0 0.03fF
C435 a_536_696# a_542_689# 0.06fF
C436 a_63_1351# a_536_696# 0.33fF
C437 a_283_1351# a_495_1121# 0.21fF
C438 c4 w_667_821# 0.03fF
C439 a_402_639# a_334_788# 0.36fF
C440 b2 a_570_1365# 0.06fF
C441 a_283_1351# a1 0.12fF
C442 a_483_781# a_542_689# 0.02fF
C443 a_530_778# w_480_1052# 0.03fF
C444 a_122_639# w_109_651# 0.03fF
C445 a_685_1058# a_720_771# 0.05fF
C446 a_678_771# gnd 0.27fF
C447 a_693_1383# a_696_771# 0.05fF
C448 w_337_1327# vdd 0.05fF
C449 a_473_1383# a_503_1351# 0.05fF
C450 a_116_696# w_221_1115# 0.06fF
C451 c0 w_480_982# 0.06fF
C452 vdd w_557_1377# 0.05fF
C453 a_381_785# w_331_1052# 0.03fF
C454 a_63_1351# a_33_1383# 0.05fF
C455 gnd a_570_1365# 0.08fF
C456 a_63_1351# a_495_1058# 0.11fF
C457 a_678_771# w_667_821# 0.10fF
C458 a_396_696# w_480_982# 0.06fF
C459 a_542_639# w_559_701# 0.06fF
C460 a_283_1351# a_256_696# 7.28fF
C461 w_117_1327# a_130_1315# 0.03fF
C462 b2 w_557_1377# 0.06fF
C463 b3 vdd 0.48fF
C464 a2 w_557_1327# 0.06fF
C465 w_18_1377# a0 0.06fF
C466 a_536_696# w_670_982# 0.06fF
C467 c0 a_116_696# 6.02fF
C468 s3 vdd 0.03fF
C469 a_685_911# a_256_696# 0.08fF
C470 a_536_696# vdd 0.85fF
C471 a_381_785# a_369_785# 0.85fF
C472 a3 vdd 0.22fF
C473 a_396_696# a_116_696# 0.41fF
C474 a_542_689# w_529_701# 0.03fF
C475 a_483_781# vdd 0.22fF
C476 w_109_701# vdd 0.05fF
C477 w_367_1377# vdd 0.11fF
C478 a_685_1121# a_503_1351# 0.21fF
C479 a_63_1351# a_256_696# 3.72fF
C480 w_109_651# vdd 0.05fF
C481 a_122_689# w_109_701# 0.03fF
C482 a_495_1121# a_518_778# 0.05fF
C483 a_63_1351# w_18_1377# 0.03fF
C484 b1 w_238_1377# 0.06fF
C485 a_495_1121# vdd 0.05fF
C486 w_147_1377# vdd 0.11fF
C487 a_744_771# a_720_771# 0.08fF
C488 a_503_1351# w_477_821# 0.06fF
C489 a_33_1383# vdd 0.05fF
C490 b3 gnd 0.21fF
C491 a_570_1365# a2 0.02fF
C492 a_495_1058# vdd 0.16fF
C493 b1 w_337_1377# 0.06fF
C494 a_253_1383# a1 0.03fF
C495 a_63_1351# a0 0.12fF
C496 vdd a1 0.22fF
C497 s3 gnd 0.13fF
C498 w_419_701# vdd 0.11fF
C499 a_696_771# a_503_1351# 0.09fF
C500 a_63_1351# a_283_1351# 0.26fF
C501 a_536_696# gnd 2.96fF
C502 s1 a_256_696# 0.12fF
C503 a3 gnd 0.76fF
C504 a_402_689# vdd 0.74fF
C505 gnd a_483_781# 0.89fF
C506 a_396_696# a_570_1365# 0.08fF
C507 a_536_696# w_670_1052# 0.06fF
C508 a_503_1351# a_542_778# 0.08fF
C509 a_483_781# w_529_651# 0.06fF
C510 b0 a_130_1365# 0.06fF
C511 w_587_1377# a_570_1365# 0.19fF
C512 w_807_1377# vdd 0.11fF
C513 a_488_778# a_503_1351# 0.54fF
C514 w_670_982# a_256_696# 0.06fF
C515 w_529_701# vdd 0.05fF
C516 a_402_639# w_389_651# 0.03fF
C517 a_570_1315# vdd 0.11fF
C518 a_350_1315# a_350_1365# 0.02fF
C519 vdd a_256_696# 1.23fF
C520 gnd a_495_1121# 0.08fF
C521 gnd a_33_1383# 0.04fF
C522 a_495_988# a_256_696# 0.17fF
C523 a_63_1351# a_259_792# 0.99fF
C524 a_495_1058# gnd 0.08fF
C525 a_262_639# s1 0.08fF
C526 gnd a1 0.76fF
C527 a_744_771# w_670_905# 0.03fF
C528 a_696_771# a_744_771# 0.08fF
C529 w_18_1377# vdd 0.14fF
C530 a_224_795# a_536_696# 0.09fF
C531 a_536_696# a_790_1315# 0.08fF
C532 a3 a_790_1315# 0.36fF
C533 s3 Gnd 1.08fF
C534 a_542_639# Gnd 1.09fF
C535 a_542_689# Gnd 0.88fF
C536 s2 Gnd 1.08fF
C537 a_402_639# Gnd 1.09fF
C538 a_402_689# Gnd 0.88fF
C539 s1 Gnd 1.08fF
C540 a_262_639# Gnd 1.09fF
C541 a_262_689# Gnd 0.88fF
C542 s0 Gnd 1.08fF
C543 a_122_639# Gnd 1.09fF
C544 a_122_689# Gnd 0.88fF
C545 c4 Gnd 2.29fF
C546 a_483_781# Gnd 3.25fF
C547 a_334_788# Gnd 3.30fF
C548 a_224_795# Gnd 3.01fF
C549 a_678_771# Gnd 0.63fF
C550 a_488_778# Gnd 0.52fF
C551 a_339_785# Gnd 0.43fF
C552 a_229_792# Gnd 0.32fF
C553 a_744_771# Gnd 1.30fF
C554 a_685_911# Gnd 0.61fF
C555 a_732_771# Gnd 2.34fF
C556 a_542_778# Gnd 2.05fF
C557 a_685_988# Gnd 0.51fF
C558 a_495_988# Gnd 0.51fF
C559 a_720_771# Gnd 3.29fF
C560 a_530_778# Gnd 2.95fF
C561 a_381_785# Gnd 2.74fF
C562 a_685_1058# Gnd 0.42fF
C563 a_495_1058# Gnd 0.42fF
C564 a_346_1058# Gnd 0.42fF
C565 a_708_771# Gnd 4.17fF
C566 a_518_778# Gnd 3.79fF
C567 a_369_785# Gnd 3.58fF
C568 a_259_792# Gnd 3.38fF
C569 a_685_1121# Gnd 0.32fF
C570 a_495_1121# Gnd 0.32fF
C571 a_346_1121# Gnd 0.32fF
C572 a_236_1121# Gnd 0.32fF
C573 c0 Gnd 18.74fF
C574 a_536_696# Gnd 21.08fF
C575 a_696_771# Gnd 15.60fF
C576 a_790_1315# Gnd 1.09fF
C577 a_693_1383# Gnd 0.32fF
C578 b3 Gnd 3.91fF
C579 a3 Gnd 3.51fF
C580 a_790_1365# Gnd 0.88fF
C581 a_396_696# Gnd 21.46fF
C582 a_503_1351# Gnd 14.24fF
C583 a_570_1315# Gnd 1.09fF
C584 a_473_1383# Gnd 0.32fF
C585 b2 Gnd 3.91fF
C586 a2 Gnd 3.51fF
C587 a_570_1365# Gnd 0.88fF
C588 a_256_696# Gnd 20.55fF
C589 a_283_1351# Gnd 13.67fF
C590 a_350_1315# Gnd 1.09fF
C591 a_253_1383# Gnd 0.32fF
C592 b1 Gnd 3.91fF
C593 a1 Gnd 3.51fF
C594 a_350_1365# Gnd 0.88fF
C595 gnd Gnd 27.15fF
C596 a_116_696# Gnd 18.02fF
C597 a_63_1351# Gnd 13.77fF
C598 vdd Gnd 24.27fF
C599 a_130_1315# Gnd 1.09fF
C600 a_33_1383# Gnd 0.32fF
C601 b0 Gnd 3.91fF
C602 a0 Gnd 3.51fF
C603 a_130_1365# Gnd 0.88fF
C604 w_529_651# Gnd 0.48fF
C605 w_389_651# Gnd 0.48fF
C606 w_249_651# Gnd 0.48fF
C607 w_109_651# Gnd 0.48fF
C608 w_559_701# Gnd 1.12fF
C609 w_529_701# Gnd 0.48fF
C610 w_419_701# Gnd 1.12fF
C611 w_389_701# Gnd 0.48fF
C612 w_279_701# Gnd 1.12fF
C613 w_249_701# Gnd 0.48fF
C614 w_139_701# Gnd 1.12fF
C615 w_109_701# Gnd 0.48fF
C616 w_667_821# Gnd 1.85fF
C617 w_477_821# Gnd 1.61fF
C618 w_328_821# Gnd 1.37fF
C619 w_218_821# Gnd 1.12fF
C620 w_670_905# Gnd 1.85fF
C621 w_670_982# Gnd 1.61fF
C622 w_480_982# Gnd 1.61fF
C623 w_670_1052# Gnd 1.37fF
C624 w_480_1052# Gnd 1.37fF
C625 w_331_1052# Gnd 1.37fF
C626 w_670_1115# Gnd 1.12fF
C627 w_480_1115# Gnd 1.12fF
C628 w_331_1115# Gnd 1.12fF
C629 w_221_1115# Gnd 1.12fF
C630 w_777_1327# Gnd 0.48fF
C631 w_557_1327# Gnd 0.48fF
C632 w_337_1327# Gnd 0.48fF
C633 w_117_1327# Gnd 0.48fF
C634 w_807_1377# Gnd 1.12fF
C635 w_777_1377# Gnd 0.48fF
C636 w_678_1377# Gnd 1.12fF
C637 w_587_1377# Gnd 1.12fF
C638 w_557_1377# Gnd 0.48fF
C639 w_458_1377# Gnd 1.12fF
C640 w_367_1377# Gnd 1.12fF
C641 w_337_1377# Gnd 0.48fF
C642 w_238_1377# Gnd 1.12fF
C643 w_147_1377# Gnd 1.12fF
C644 w_117_1377# Gnd 0.48fF
C645 w_18_1377# Gnd 1.12fF

** Analysis **
.tran 1p 80n

** Plotting **
.control
set hcopypscolor=1
set color0=white
set color1=black
run
set curplottitle="2020102037"
plot a0 a1+2 a2+4 a3+6
plot b0 b1+2 b2+4 b3+6
plot s0 s1+2 s2+4 s3+6 c4+8
.endc

.end