magic
tech scmos
timestamp 1638582313
<< nwell >>
rect 0 0 56 20
<< ntransistor >>
rect 13 -26 15 -22
rect 25 -26 27 -22
rect 43 -26 45 -22
<< ptransistor >>
rect 13 6 15 14
rect 25 6 27 14
rect 43 6 45 14
<< ndiffusion >>
rect 10 -26 13 -22
rect 15 -26 25 -22
rect 27 -26 30 -22
rect 42 -26 43 -22
rect 45 -26 46 -22
<< pdiffusion >>
rect 10 6 13 14
rect 15 6 18 14
rect 22 6 25 14
rect 27 6 30 14
rect 42 6 43 14
rect 45 6 46 14
<< ndcontact >>
rect 6 -26 10 -22
rect 30 -26 34 -22
rect 38 -26 42 -22
rect 46 -26 50 -22
<< pdcontact >>
rect 6 6 10 14
rect 18 6 22 14
rect 30 6 34 14
rect 38 6 42 14
rect 46 6 50 14
<< polysilicon >>
rect 13 14 15 17
rect 25 14 27 17
rect 43 14 45 17
rect 13 -22 15 6
rect 25 -22 27 6
rect 43 -22 45 6
rect 13 -29 15 -26
rect 25 -29 27 -26
rect 43 -29 45 -26
<< polycontact >>
rect 9 -5 13 -1
rect 21 -12 25 -8
rect 39 -13 43 -9
<< metal1 >>
rect 0 20 56 24
rect 6 14 10 20
rect 30 14 34 20
rect 38 14 42 20
rect 18 -1 22 6
rect 0 -5 9 -1
rect 18 -5 34 -1
rect 0 -12 21 -8
rect 30 -9 34 -5
rect 46 -9 50 6
rect 30 -13 39 -9
rect 46 -13 56 -9
rect 30 -22 34 -13
rect 46 -22 50 -13
rect 6 -30 10 -26
rect 38 -30 42 -26
rect 0 -34 56 -30
<< labels >>
rlabel metal1 0 -5 4 -1 3 in1
rlabel metal1 0 -12 4 -8 3 in2
rlabel metal1 0 20 56 24 5 vdd
rlabel metal1 52 -13 56 -9 7 out
rlabel metal1 0 -34 56 -30 1 gnd
<< end >>
