* SPICE3 file created from or2.ext - technology: scmos

.option scale=0.09u

M1000 a_15_6# in1 vdd w_0_0# pfet w=8 l=2
+  ad=80 pd=36 as=96 ps=56
M1001 a_15_n26# in2 a_15_6# w_0_0# pfet w=8 l=2
+  ad=56 pd=30 as=0 ps=0
M1002 a_15_n26# in1 gnd Gnd nfet w=4 l=2
+  ad=40 pd=28 as=76 ps=62
M1003 out a_15_n26# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1004 out a_15_n26# vdd w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1005 gnd in2 a_15_n26# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out vdd 0.11fF
C1 a_15_n26# in2 0.21fF
C2 a_15_n26# vdd 0.11fF
C3 w_0_0# in2 0.06fF
C4 w_0_0# vdd 0.11fF
C5 w_0_0# in1 0.06fF
C6 in1 in2 0.27fF
C7 in1 vdd 0.02fF
C8 a_15_n26# out 0.05fF
C9 w_0_0# out 0.03fF
C10 out gnd 0.08fF
C11 w_0_0# a_15_n26# 0.10fF
C12 a_15_n26# gnd 0.10fF
C13 gnd Gnd 0.24fF
C14 out Gnd 0.10fF
C15 vdd Gnd 0.13fF
C16 a_15_n26# Gnd 0.32fF
C17 in2 Gnd 0.26fF
C18 in1 Gnd 0.23fF
C19 w_0_0# Gnd 1.12fF
