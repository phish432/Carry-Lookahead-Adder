magic
tech scmos
timestamp 1638840513
<< nwell >>
rect 139 86 163 106
rect 169 86 225 106
rect 279 86 303 106
rect 309 86 365 106
rect 419 86 443 106
rect 449 86 505 106
rect 559 86 583 106
rect 589 86 645 106
rect 139 36 163 56
rect 279 36 303 56
rect 419 36 443 56
rect 559 36 583 56
<< ntransistor >>
rect 150 74 152 78
rect 290 74 292 78
rect 430 74 432 78
rect 570 74 572 78
rect 150 24 152 28
rect 181 24 183 28
rect 191 24 193 28
rect 201 24 203 28
rect 211 24 213 28
rect 290 24 292 28
rect 321 24 323 28
rect 331 24 333 28
rect 341 24 343 28
rect 351 24 353 28
rect 430 24 432 28
rect 461 24 463 28
rect 471 24 473 28
rect 481 24 483 28
rect 491 24 493 28
rect 570 24 572 28
rect 601 24 603 28
rect 611 24 613 28
rect 621 24 623 28
rect 631 24 633 28
<< ptransistor >>
rect 150 92 152 100
rect 181 92 183 100
rect 191 92 193 100
rect 201 92 203 100
rect 211 92 213 100
rect 150 42 152 50
rect 290 92 292 100
rect 321 92 323 100
rect 331 92 333 100
rect 341 92 343 100
rect 351 92 353 100
rect 290 42 292 50
rect 430 92 432 100
rect 461 92 463 100
rect 471 92 473 100
rect 481 92 483 100
rect 491 92 493 100
rect 430 42 432 50
rect 570 92 572 100
rect 601 92 603 100
rect 611 92 613 100
rect 621 92 623 100
rect 631 92 633 100
rect 570 42 572 50
<< ndiffusion >>
rect 149 74 150 78
rect 152 74 153 78
rect 289 74 290 78
rect 292 74 293 78
rect 429 74 430 78
rect 432 74 433 78
rect 569 74 570 78
rect 572 74 573 78
rect 149 24 150 28
rect 152 24 153 28
rect 179 24 181 28
rect 183 24 191 28
rect 193 24 195 28
rect 199 24 201 28
rect 203 24 211 28
rect 213 24 215 28
rect 289 24 290 28
rect 292 24 293 28
rect 319 24 321 28
rect 323 24 331 28
rect 333 24 335 28
rect 339 24 341 28
rect 343 24 351 28
rect 353 24 355 28
rect 429 24 430 28
rect 432 24 433 28
rect 459 24 461 28
rect 463 24 471 28
rect 473 24 475 28
rect 479 24 481 28
rect 483 24 491 28
rect 493 24 495 28
rect 569 24 570 28
rect 572 24 573 28
rect 599 24 601 28
rect 603 24 611 28
rect 613 24 615 28
rect 619 24 621 28
rect 623 24 631 28
rect 633 24 635 28
<< pdiffusion >>
rect 149 92 150 100
rect 152 92 153 100
rect 179 92 181 100
rect 183 92 191 100
rect 193 92 195 100
rect 199 92 201 100
rect 203 92 211 100
rect 213 92 215 100
rect 149 42 150 50
rect 152 42 153 50
rect 289 92 290 100
rect 292 92 293 100
rect 319 92 321 100
rect 323 92 331 100
rect 333 92 335 100
rect 339 92 341 100
rect 343 92 351 100
rect 353 92 355 100
rect 289 42 290 50
rect 292 42 293 50
rect 429 92 430 100
rect 432 92 433 100
rect 459 92 461 100
rect 463 92 471 100
rect 473 92 475 100
rect 479 92 481 100
rect 483 92 491 100
rect 493 92 495 100
rect 429 42 430 50
rect 432 42 433 50
rect 569 92 570 100
rect 572 92 573 100
rect 599 92 601 100
rect 603 92 611 100
rect 613 92 615 100
rect 619 92 621 100
rect 623 92 631 100
rect 633 92 635 100
rect 569 42 570 50
rect 572 42 573 50
<< ndcontact >>
rect 145 74 149 78
rect 153 74 157 78
rect 285 74 289 78
rect 293 74 297 78
rect 425 74 429 78
rect 433 74 437 78
rect 565 74 569 78
rect 573 74 577 78
rect 145 24 149 28
rect 153 24 157 28
rect 175 24 179 28
rect 195 24 199 28
rect 215 24 219 28
rect 285 24 289 28
rect 293 24 297 28
rect 315 24 319 28
rect 335 24 339 28
rect 355 24 359 28
rect 425 24 429 28
rect 433 24 437 28
rect 455 24 459 28
rect 475 24 479 28
rect 495 24 499 28
rect 565 24 569 28
rect 573 24 577 28
rect 595 24 599 28
rect 615 24 619 28
rect 635 24 639 28
<< pdcontact >>
rect 145 92 149 100
rect 153 92 157 100
rect 175 92 179 100
rect 195 92 199 100
rect 215 92 219 100
rect 145 42 149 50
rect 153 42 157 50
rect 285 92 289 100
rect 293 92 297 100
rect 315 92 319 100
rect 335 92 339 100
rect 355 92 359 100
rect 285 42 289 50
rect 293 42 297 50
rect 425 92 429 100
rect 433 92 437 100
rect 455 92 459 100
rect 475 92 479 100
rect 495 92 499 100
rect 425 42 429 50
rect 433 42 437 50
rect 565 92 569 100
rect 573 92 577 100
rect 595 92 599 100
rect 615 92 619 100
rect 635 92 639 100
rect 565 42 569 50
rect 573 42 577 50
<< polysilicon >>
rect 181 110 223 112
rect 150 100 152 103
rect 181 100 183 110
rect 191 100 193 103
rect 201 100 203 103
rect 211 100 213 103
rect 150 78 152 92
rect 181 81 183 92
rect 191 77 193 92
rect 181 75 193 77
rect 150 71 152 74
rect 150 50 152 53
rect 150 28 152 42
rect 181 28 183 75
rect 201 72 203 92
rect 191 70 203 72
rect 191 28 193 70
rect 211 38 213 92
rect 201 36 213 38
rect 201 28 203 36
rect 221 33 223 110
rect 321 110 363 112
rect 290 100 292 103
rect 321 100 323 110
rect 331 100 333 103
rect 341 100 343 103
rect 351 100 353 103
rect 290 78 292 92
rect 321 81 323 92
rect 331 77 333 92
rect 321 75 333 77
rect 290 71 292 74
rect 290 50 292 53
rect 211 31 223 33
rect 211 28 213 31
rect 290 28 292 42
rect 321 28 323 75
rect 341 72 343 92
rect 331 70 343 72
rect 331 28 333 70
rect 351 38 353 92
rect 341 36 353 38
rect 341 28 343 36
rect 361 33 363 110
rect 461 110 503 112
rect 430 100 432 103
rect 461 100 463 110
rect 471 100 473 103
rect 481 100 483 103
rect 491 100 493 103
rect 430 78 432 92
rect 461 81 463 92
rect 471 77 473 92
rect 461 75 473 77
rect 430 71 432 74
rect 430 50 432 53
rect 351 31 363 33
rect 351 28 353 31
rect 430 28 432 42
rect 461 28 463 75
rect 481 72 483 92
rect 471 70 483 72
rect 471 28 473 70
rect 491 38 493 92
rect 481 36 493 38
rect 481 28 483 36
rect 501 33 503 110
rect 601 110 643 112
rect 570 100 572 103
rect 601 100 603 110
rect 611 100 613 103
rect 621 100 623 103
rect 631 100 633 103
rect 570 78 572 92
rect 601 81 603 92
rect 611 77 613 92
rect 601 75 613 77
rect 570 71 572 74
rect 570 50 572 53
rect 491 31 503 33
rect 491 28 493 31
rect 570 28 572 42
rect 601 28 603 75
rect 621 72 623 92
rect 611 70 623 72
rect 611 28 613 70
rect 631 38 633 92
rect 621 36 633 38
rect 621 28 623 36
rect 641 33 643 110
rect 631 31 643 33
rect 631 28 633 31
rect 150 21 152 24
rect 181 8 183 24
rect 191 21 193 24
rect 201 0 203 24
rect 211 21 213 24
rect 290 21 292 24
rect 321 8 323 24
rect 331 21 333 24
rect 341 0 343 24
rect 351 21 353 24
rect 430 21 432 24
rect 461 8 463 24
rect 471 21 473 24
rect 481 0 483 24
rect 491 21 493 24
rect 570 21 572 24
rect 601 8 603 24
rect 611 21 613 24
rect 621 0 623 24
rect 631 21 633 24
<< polycontact >>
rect 146 81 150 85
rect 177 81 181 85
rect 146 31 150 35
rect 187 61 191 65
rect 286 81 290 85
rect 317 81 321 85
rect 286 31 290 35
rect 327 61 331 65
rect 426 81 430 85
rect 457 81 461 85
rect 426 31 430 35
rect 467 61 471 65
rect 566 81 570 85
rect 597 81 601 85
rect 566 31 570 35
rect 607 61 611 65
rect 177 8 181 12
rect 197 0 201 4
rect 317 8 321 12
rect 337 0 341 4
rect 457 8 461 12
rect 477 0 481 4
rect 597 8 601 12
rect 617 0 621 4
<< metal1 >>
rect 116 106 645 110
rect 116 81 120 85
rect 130 60 134 106
rect 145 100 149 106
rect 175 100 179 106
rect 215 100 219 106
rect 153 85 157 92
rect 142 81 146 85
rect 153 81 177 85
rect 153 78 157 81
rect 145 70 149 74
rect 139 66 172 70
rect 130 56 163 60
rect 145 50 149 56
rect 153 35 157 42
rect 108 31 129 35
rect 134 31 146 35
rect 153 31 160 35
rect 153 28 157 31
rect 145 20 149 24
rect 168 20 172 66
rect 180 61 187 65
rect 195 59 199 92
rect 256 81 260 85
rect 270 60 274 106
rect 285 100 289 106
rect 315 100 319 106
rect 355 100 359 106
rect 293 85 297 92
rect 282 81 286 85
rect 293 81 317 85
rect 293 78 297 81
rect 285 70 289 74
rect 279 66 312 70
rect 195 55 227 59
rect 195 28 199 55
rect 270 56 303 60
rect 285 50 289 56
rect 293 35 297 42
rect 248 31 269 35
rect 274 31 286 35
rect 293 31 300 35
rect 293 28 297 31
rect 175 20 179 24
rect 215 20 219 24
rect 285 20 289 24
rect 308 20 312 66
rect 320 61 327 65
rect 335 59 339 92
rect 396 81 400 85
rect 410 60 414 106
rect 425 100 429 106
rect 455 100 459 106
rect 495 100 499 106
rect 433 85 437 92
rect 422 81 426 85
rect 433 81 457 85
rect 433 78 437 81
rect 425 70 429 74
rect 419 66 452 70
rect 335 55 367 59
rect 335 28 339 55
rect 410 56 443 60
rect 425 50 429 56
rect 433 35 437 42
rect 388 31 409 35
rect 414 31 426 35
rect 433 31 440 35
rect 433 28 437 31
rect 315 20 319 24
rect 355 20 359 24
rect 425 20 429 24
rect 448 20 452 66
rect 460 61 467 65
rect 475 59 479 92
rect 536 81 540 85
rect 550 60 554 106
rect 565 100 569 106
rect 595 100 599 106
rect 635 100 639 106
rect 573 85 577 92
rect 562 81 566 85
rect 573 81 597 85
rect 573 78 577 81
rect 565 70 569 74
rect 559 66 592 70
rect 475 55 507 59
rect 475 28 479 55
rect 550 56 583 60
rect 565 50 569 56
rect 573 35 577 42
rect 528 31 549 35
rect 554 31 566 35
rect 573 31 580 35
rect 573 28 577 31
rect 455 20 459 24
rect 495 20 499 24
rect 565 20 569 24
rect 588 20 592 66
rect 600 61 607 65
rect 615 59 619 92
rect 615 55 647 59
rect 615 28 619 55
rect 595 20 599 24
rect 635 20 639 24
rect 116 16 645 20
rect 135 8 177 12
rect 275 8 317 12
rect 415 8 457 12
rect 555 8 597 12
rect 166 0 197 4
rect 306 0 337 4
rect 446 0 477 4
rect 586 0 617 4
<< m2contact >>
rect 111 81 116 86
rect 120 80 125 85
rect 137 80 142 85
rect 103 31 108 36
rect 129 30 134 35
rect 160 30 165 35
rect 175 60 180 65
rect 251 81 256 86
rect 260 80 265 85
rect 277 80 282 85
rect 227 54 232 59
rect 243 31 248 36
rect 269 30 274 35
rect 300 30 305 35
rect 315 60 320 65
rect 391 81 396 86
rect 400 80 405 85
rect 417 80 422 85
rect 367 54 372 59
rect 383 31 388 36
rect 409 30 414 35
rect 440 30 445 35
rect 455 60 460 65
rect 531 81 536 86
rect 540 80 545 85
rect 557 80 562 85
rect 507 54 512 59
rect 523 31 528 36
rect 549 30 554 35
rect 580 30 585 35
rect 595 60 600 65
rect 647 54 652 59
rect 130 8 135 13
rect 270 8 275 13
rect 410 8 415 13
rect 550 8 555 13
rect 161 0 166 5
rect 301 0 306 5
rect 441 0 446 5
rect 581 0 586 5
<< metal2 >>
rect 103 36 107 124
rect 111 86 115 124
rect 125 80 137 84
rect 121 65 125 80
rect 121 61 175 65
rect 130 13 134 30
rect 161 5 165 30
rect 228 -8 232 54
rect 243 36 247 124
rect 251 86 255 124
rect 265 80 277 84
rect 261 65 265 80
rect 261 61 315 65
rect 270 13 274 30
rect 301 5 305 30
rect 368 -14 372 54
rect 383 36 387 124
rect 391 86 395 124
rect 405 80 417 84
rect 401 65 405 80
rect 401 61 455 65
rect 410 13 414 30
rect 441 5 445 30
rect 508 -14 512 54
rect 523 36 527 124
rect 531 86 535 124
rect 545 80 557 84
rect 541 65 545 80
rect 541 61 595 65
rect 550 13 554 30
rect 581 5 585 30
rect 648 -14 652 54
<< labels >>
rlabel metal2 243 120 247 124 5 p1
rlabel metal2 251 120 255 124 5 c1
rlabel metal2 383 120 387 124 5 p2
rlabel metal2 391 120 395 124 5 c2
rlabel metal2 523 120 527 124 5 p3
rlabel metal2 531 120 535 124 5 c3
rlabel metal2 648 -14 652 -10 8 s3
rlabel metal2 508 -14 512 -10 1 s2
rlabel metal2 368 -14 372 -10 1 s1
rlabel metal1 116 106 645 110 1 vdd
rlabel metal1 116 16 645 20 1 gnd
rlabel metal2 103 120 107 124 4 p0
rlabel metal2 111 120 115 124 5 c0
rlabel metal2 228 -8 232 -4 1 s0
<< end >>
